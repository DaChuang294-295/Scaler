library verilog;
use verilog.vl_types.all;
entity OSC is
    port(
        outclk          : out    vl_logic
    );
end OSC;
