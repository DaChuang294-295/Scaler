library verilog;
use verilog.vl_types.all;
entity GND is
    port(
        Y               : out    vl_logic
    );
end GND;
