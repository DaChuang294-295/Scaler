library verilog;
use verilog.vl_types.all;
entity emb_16_2k is
    port(
        clka            : in     vl_logic;
        cea             : in     vl_logic;
        wea             : in     vl_logic;
        aa              : in     vl_logic_vector(10 downto 0);
        da              : in     vl_logic_vector(15 downto 0);
        qa              : out    vl_logic_vector(15 downto 0);
        clkb            : in     vl_logic;
        ceb             : in     vl_logic;
        web             : in     vl_logic;
        ab              : in     vl_logic_vector(10 downto 0);
        db              : in     vl_logic_vector(15 downto 0);
        qb              : out    vl_logic_vector(15 downto 0)
    );
end emb_16_2k;
