library verilog;
use verilog.vl_types.all;
entity gbuf_v1_1 is
    port(
        I               : in     vl_logic;
        O               : out    vl_logic
    );
end gbuf_v1_1;
