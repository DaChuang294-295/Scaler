library verilog;
use verilog.vl_types.all;
entity m7s_hm2pm_if_async is
    generic(
        IDLE            : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        BUSY            : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        NONSEQ          : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        SEQ             : vl_logic_vector(0 to 1) := (Hi1, Hi1);
        SINGLE          : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        INCR            : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        WRAP4           : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        INCR4           : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        WRAP8           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        INCR8           : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        WRAP16          : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        INCR16          : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        H_IDLE          : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        H_RDATA         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        H_WDATA         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        H_WDATA_WAIT    : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        P_IDLE          : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        P_CMD           : vl_logic_vector(0 to 1) := (Hi0, Hi1);
        P_WDATA         : vl_logic_vector(0 to 1) := (Hi1, Hi0);
        P_RDATA         : vl_logic_vector(0 to 1) := (Hi1, Hi1)
    );
    port(
        clk_pbus        : in     vl_logic;
        rst_pbus_n      : in     vl_logic;
        clk_ahb         : in     vl_logic;
        rst_ahb_n       : in     vl_logic;
        ahb_mastlock    : in     vl_logic;
        ahb_prot        : in     vl_logic_vector(3 downto 0);
        ahb_size        : in     vl_logic_vector(2 downto 0);
        ahb_addr        : in     vl_logic_vector(31 downto 0);
        ahb_write       : in     vl_logic;
        ahb_burst       : in     vl_logic_vector(2 downto 0);
        ahb_trans       : in     vl_logic_vector(1 downto 0);
        ahb_wdata       : in     vl_logic_vector(31 downto 0);
        ahb_ready       : out    vl_logic;
        ahb_resp        : out    vl_logic;
        ahb_rdata       : out    vl_logic_vector(31 downto 0);
        pbus_aid        : out    vl_logic_vector(3 downto 0);
        pbus_addr       : out    vl_logic_vector(31 downto 0);
        pbus_write      : out    vl_logic;
        pbus_length     : out    vl_logic_vector(3 downto 0);
        pbus_wbyte_en   : out    vl_logic_vector(3 downto 0);
        pbus_type_burst : out    vl_logic_vector(1 downto 0);
        pbus_avalid     : out    vl_logic;
        pbus_aready     : in     vl_logic;
        pbus_wdata      : out    vl_logic_vector(31 downto 0);
        pbus_wvalid     : out    vl_logic;
        pbus_wready     : in     vl_logic;
        pbus_did        : in     vl_logic_vector(3 downto 0);
        pbus_rdata      : in     vl_logic_vector(31 downto 0);
        pbus_rready     : out    vl_logic;
        pbus_rvalid     : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of BUSY : constant is 1;
    attribute mti_svvh_generic_type of NONSEQ : constant is 1;
    attribute mti_svvh_generic_type of SEQ : constant is 1;
    attribute mti_svvh_generic_type of SINGLE : constant is 1;
    attribute mti_svvh_generic_type of INCR : constant is 1;
    attribute mti_svvh_generic_type of WRAP4 : constant is 1;
    attribute mti_svvh_generic_type of INCR4 : constant is 1;
    attribute mti_svvh_generic_type of WRAP8 : constant is 1;
    attribute mti_svvh_generic_type of INCR8 : constant is 1;
    attribute mti_svvh_generic_type of WRAP16 : constant is 1;
    attribute mti_svvh_generic_type of INCR16 : constant is 1;
    attribute mti_svvh_generic_type of H_IDLE : constant is 1;
    attribute mti_svvh_generic_type of H_RDATA : constant is 1;
    attribute mti_svvh_generic_type of H_WDATA : constant is 1;
    attribute mti_svvh_generic_type of H_WDATA_WAIT : constant is 1;
    attribute mti_svvh_generic_type of P_IDLE : constant is 1;
    attribute mti_svvh_generic_type of P_CMD : constant is 1;
    attribute mti_svvh_generic_type of P_WDATA : constant is 1;
    attribute mti_svvh_generic_type of P_RDATA : constant is 1;
end m7s_hm2pm_if_async;
