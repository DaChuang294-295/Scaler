library verilog;
use verilog.vl_types.all;
entity por_v1_1 is
    port(
        O               : out    vl_logic
    );
end por_v1_1;
