library verilog;
use verilog.vl_types.all;
entity GBUF is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end GBUF;
