library verilog;
use verilog.vl_types.all;
entity M7S_SOC is
    generic(
        SIM_FIFO        : integer := 0;
        START_ADDR      : vl_logic_vector(31 downto 0) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        use_arm         : vl_logic := Hi1;
        use_clk_arm     : vl_logic := Hi1;
        use_pbus0       : vl_logic := Hi1;
        use_pbus1       : vl_logic := Hi1;
        use_on_chip_eth : vl_logic := Hi0;
        use_on_chip_usb : vl_logic := Hi0;
        use_on_chip_ddr_ctrl: vl_logic := Hi0;
        use_on_chip_adc : vl_logic_vector(0 to 11) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        use_uart_io     : vl_logic := Hi0;
        use_arm_nmi     : vl_logic := Hi0;
        on_chip_ddr_ctrl_mode: string  := "";
        on_chip_eth_mode: string  := "";
        program_file    : string  := ""
    );
    port(
        fp2soc_rst_n    : in     vl_logic;
        c2r1_dll_clk    : in     vl_logic;
        fp_lvds_sclk    : in     vl_logic;
        fp_clk_sys      : in     vl_logic;
        fp_clk_adc      : in     vl_logic;
        fp_clk_arm      : in     vl_logic;
        fp_clk_usb      : in     vl_logic;
        clk_eth_tx      : in     vl_logic;
        gpio_0_out_o    : out    vl_logic_vector(31 downto 0);
        gpio_0_oe_o     : out    vl_logic_vector(31 downto 0);
        gpio_0_in_i     : in     vl_logic_vector(31 downto 0);
        i2c0_scl_oe_o   : out    vl_logic;
        i2c0_sda_oe_o   : out    vl_logic;
        i2c0_scl_i      : in     vl_logic;
        i2c0_sda_i      : in     vl_logic;
        i2c1_scl_oe_o   : out    vl_logic;
        i2c1_sda_oe_o   : out    vl_logic;
        i2c1_scl_i      : in     vl_logic;
        i2c1_sda_i      : in     vl_logic;
        uart0_rts_o     : out    vl_logic;
        uart0_txd_o     : out    vl_logic;
        uart0_cts_i     : in     vl_logic;
        uart0_rxd_i     : in     vl_logic;
        uart1_rts_o     : out    vl_logic;
        uart1_txd_o     : out    vl_logic;
        uart1_cts_i     : in     vl_logic;
        uart1_rxd_i     : in     vl_logic;
        spi0_mosi       : out    vl_logic;
        spi0_sck        : out    vl_logic;
        spi0_ssn        : out    vl_logic;
        spi0_miso       : in     vl_logic;
        spi1_mosi       : out    vl_logic;
        spi1_sck        : out    vl_logic;
        spi1_ssn        : out    vl_logic;
        spi1_miso       : in     vl_logic;
        pad_can0_o_clk  : out    vl_logic;
        pad_can0_o_tx1  : out    vl_logic;
        pad_can0_o_tx0  : out    vl_logic;
        pad_can0_oen_tx1: out    vl_logic;
        pad_can0_oen_tx0: out    vl_logic;
        pad_can0_i_rx0  : in     vl_logic;
        pad_can1_o_clk  : out    vl_logic;
        pad_can1_o_tx1  : out    vl_logic;
        pad_can1_o_tx0  : out    vl_logic;
        pad_can1_oen_tx1: out    vl_logic;
        pad_can1_oen_tx0: out    vl_logic;
        pad_can1_i_rx0  : in     vl_logic;
        clk_ahb_fp1     : in     vl_logic;
        rst_ahb_fp1_n   : in     vl_logic;
        fp1_m_ahb_mastlock: in     vl_logic;
        fp1_m_ahb_prot  : in     vl_logic_vector(3 downto 0);
        fp1_m_ahb_size  : in     vl_logic_vector(2 downto 0);
        fp1_m_ahb_addr  : in     vl_logic_vector(31 downto 0);
        fp1_m_ahb_write : in     vl_logic;
        fp1_m_ahb_burst : in     vl_logic_vector(2 downto 0);
        fp1_m_ahb_trans : in     vl_logic_vector(1 downto 0);
        fp1_m_ahb_wdata : in     vl_logic_vector(31 downto 0);
        fp1_m_ahb_ready : out    vl_logic;
        fp1_m_ahb_resp  : out    vl_logic;
        fp1_m_ahb_rdata : out    vl_logic_vector(31 downto 0);
        fp1_s_ahb_mastlock: out    vl_logic;
        fp1_s_ahb_prot  : out    vl_logic_vector(3 downto 0);
        fp1_s_ahb_size  : out    vl_logic_vector(2 downto 0);
        fp1_s_ahb_sel   : out    vl_logic;
        fp1_s_ahb_addr  : out    vl_logic_vector(31 downto 0);
        fp1_s_ahb_write : out    vl_logic;
        fp1_s_ahb_burst : out    vl_logic_vector(2 downto 0);
        fp1_s_ahb_trans : out    vl_logic_vector(1 downto 0);
        fp1_s_ahb_wdata : out    vl_logic_vector(31 downto 0);
        fp1_s_ahb_readyout: in     vl_logic;
        fp1_s_ahb_resp  : in     vl_logic;
        fp1_s_ahb_rdata : in     vl_logic_vector(31 downto 0);
        clk_ahb_fp0     : in     vl_logic;
        rst_ahb_fp0_n   : in     vl_logic;
        fp0_m_ahb_mastlock: in     vl_logic;
        fp0_m_ahb_prot  : in     vl_logic_vector(3 downto 0);
        fp0_m_ahb_size  : in     vl_logic_vector(2 downto 0);
        fp0_m_ahb_addr  : in     vl_logic_vector(31 downto 0);
        fp0_m_ahb_write : in     vl_logic;
        fp0_m_ahb_burst : in     vl_logic_vector(2 downto 0);
        fp0_m_ahb_trans : in     vl_logic_vector(1 downto 0);
        fp0_m_ahb_wdata : in     vl_logic_vector(31 downto 0);
        fp0_m_ahb_ready : out    vl_logic;
        fp0_m_ahb_resp  : out    vl_logic;
        fp0_m_ahb_rdata : out    vl_logic_vector(31 downto 0);
        fp0_s_ahb_mastlock: out    vl_logic;
        fp0_s_ahb_prot  : out    vl_logic_vector(3 downto 0);
        fp0_s_ahb_size  : out    vl_logic_vector(2 downto 0);
        fp0_s_ahb_sel   : out    vl_logic;
        fp0_s_ahb_addr  : out    vl_logic_vector(31 downto 0);
        fp0_s_ahb_write : out    vl_logic;
        fp0_s_ahb_burst : out    vl_logic_vector(2 downto 0);
        fp0_s_ahb_trans : out    vl_logic_vector(1 downto 0);
        fp0_s_ahb_wdata : out    vl_logic_vector(31 downto 0);
        fp0_s_ahb_readyout: in     vl_logic;
        fp0_s_ahb_resp  : in     vl_logic;
        fp0_s_ahb_rdata : in     vl_logic_vector(31 downto 0);
        fp_INTNMI       : in     vl_logic_vector(15 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SIM_FIFO : constant is 1;
    attribute mti_svvh_generic_type of START_ADDR : constant is 1;
    attribute mti_svvh_generic_type of use_arm : constant is 1;
    attribute mti_svvh_generic_type of use_clk_arm : constant is 1;
    attribute mti_svvh_generic_type of use_pbus0 : constant is 1;
    attribute mti_svvh_generic_type of use_pbus1 : constant is 1;
    attribute mti_svvh_generic_type of use_on_chip_eth : constant is 1;
    attribute mti_svvh_generic_type of use_on_chip_usb : constant is 1;
    attribute mti_svvh_generic_type of use_on_chip_ddr_ctrl : constant is 1;
    attribute mti_svvh_generic_type of use_on_chip_adc : constant is 1;
    attribute mti_svvh_generic_type of use_uart_io : constant is 1;
    attribute mti_svvh_generic_type of use_arm_nmi : constant is 1;
    attribute mti_svvh_generic_type of on_chip_ddr_ctrl_mode : constant is 1;
    attribute mti_svvh_generic_type of on_chip_eth_mode : constant is 1;
    attribute mti_svvh_generic_type of program_file : constant is 1;
end M7S_SOC;
