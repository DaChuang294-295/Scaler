library verilog;
use verilog.vl_types.all;
entity M7S_POR is
    port(
        z0              : out    vl_logic
    );
end M7S_POR;
