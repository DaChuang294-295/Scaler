library verilog;
use verilog.vl_types.all;
entity M7S_IO_PCISG is
    generic(
        cfg_nc          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ns_lv_fastestn  : vl_logic := Hi0;
        cfg_userio_en   : vl_logic := Hi0;
        ns_lv_cfg       : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pdr_cfg         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ndr_cfg         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        keep_cfg        : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        rx_dig_en_cfg   : vl_logic := Hi0;
        in_del          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        out_del         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        vpci_en         : vl_logic := Hi0;
        cfg_oen_inv     : vl_logic := Hi0;
        cfg_oen_sel     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_od_inv      : vl_logic := Hi0;
        cfg_od_sel      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_id_sel      : vl_logic := Hi0;
        cfg_fclk_inv    : vl_logic := Hi0;
        cfg_fclk_gate_sel: vl_logic := Hi0;
        cfg_fclk_en     : vl_logic := Hi0;
        cfg_rstn_inv    : vl_logic := Hi0;
        cfg_oen_rstn_en : vl_logic := Hi0;
        cfg_od_rstn_en  : vl_logic := Hi0;
        cfg_id_rstn_en  : vl_logic := Hi0;
        cfg_setn_inv    : vl_logic := Hi0;
        cfg_oen_setn_en : vl_logic := Hi0;
        cfg_od_setn_en  : vl_logic := Hi0;
        cfg_id_setn_en  : vl_logic := Hi0;
        optional_function: string  := ""
    );
    port(
        id              : out    vl_logic;
        clk             : in     vl_logic;
        clk_en          : in     vl_logic;
        rstn            : in     vl_logic;
        setn            : in     vl_logic;
        od              : in     vl_logic;
        oen             : in     vl_logic;
        PAD             : inout  vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of cfg_nc : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_fastestn : constant is 1;
    attribute mti_svvh_generic_type of cfg_userio_en : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_cfg : constant is 1;
    attribute mti_svvh_generic_type of pdr_cfg : constant is 1;
    attribute mti_svvh_generic_type of ndr_cfg : constant is 1;
    attribute mti_svvh_generic_type of keep_cfg : constant is 1;
    attribute mti_svvh_generic_type of rx_dig_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of in_del : constant is 1;
    attribute mti_svvh_generic_type of out_del : constant is 1;
    attribute mti_svvh_generic_type of vpci_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_gate_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_rstn_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_setn_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_setn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_setn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_setn_en : constant is 1;
    attribute mti_svvh_generic_type of optional_function : constant is 1;
end M7S_IO_PCISG;
