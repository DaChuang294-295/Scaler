library verilog;
use verilog.vl_types.all;
entity PLL_SIM is
    generic(
        MAX_INPUT_PERIOD: integer := 500;
        MIN_INPUT_PERIOD: integer := 2;
        MAX_PFD_PERIOD  : integer := 500;
        MIN_PFD_PERIOD  : real    := 2.500000;
        MAX_VCO_PERIOD  : real    := 1.667000;
        MIN_VCO_PERIOD  : real    := 0.800000;
        MAX_OUTPUT_PERIOD: integer := 100;
        MIN_OUTPUT_PERIOD: real    := 0.800000;
        LOCK_TIME       : integer := 20
    );
    port(
        VDDIO           : in     vl_logic;
        VSSIO           : in     vl_logic;
        DVDD            : in     vl_logic;
        DVSS            : in     vl_logic;
        AVSS_VCO        : in     vl_logic;
        AVSS            : in     vl_logic;
        PLLCK0          : in     vl_logic;
        PLLCK1          : in     vl_logic;
        CFBCK           : in     vl_logic;
        VREF            : in     vl_logic;
        CO0             : out    vl_logic;
        CO1             : out    vl_logic;
        CO2             : out    vl_logic;
        CO3             : out    vl_logic;
        PLOCK           : out    vl_logic;
        ACTIVECK        : out    vl_logic;
        ATEST_PLL       : out    vl_logic;
        DTEST_PLL       : out    vl_logic;
        PDB             : in     vl_logic;
        RSTPLL          : in     vl_logic;
        MKEN0           : in     vl_logic;
        MKEN1           : in     vl_logic;
        MKEN2           : in     vl_logic;
        MKEN3           : in     vl_logic;
        BPS0            : in     vl_logic;
        BPS1            : in     vl_logic;
        BPS2            : in     vl_logic;
        BPS3            : in     vl_logic;
        DIVN            : in     vl_logic_vector(7 downto 0);
        DIVM            : in     vl_logic_vector(7 downto 0);
        DIVC0           : in     vl_logic_vector(7 downto 0);
        DIVC1           : in     vl_logic_vector(7 downto 0);
        DIVC2           : in     vl_logic_vector(7 downto 0);
        DIVC3           : in     vl_logic_vector(7 downto 0);
        CO0DLY          : in     vl_logic_vector(7 downto 0);
        CO1DLY          : in     vl_logic_vector(7 downto 0);
        CO2DLY          : in     vl_logic_vector(7 downto 0);
        CO3DLY          : in     vl_logic_vector(7 downto 0);
        SEL_FBPATH      : in     vl_logic;
        DIVMP           : in     vl_logic_vector(2 downto 0);
        SEL_C0PHASE     : in     vl_logic_vector(2 downto 0);
        SEL_C1PHASE     : in     vl_logic_vector(2 downto 0);
        SEL_C2PHASE     : in     vl_logic_vector(2 downto 0);
        SEL_C3PHASE     : in     vl_logic_vector(2 downto 0);
        MP_AUTOR_EN     : in     vl_logic;
        LPF             : in     vl_logic_vector(1 downto 0);
        VRSEL           : in     vl_logic_vector(1 downto 0);
        CPSEL_CR        : in     vl_logic_vector(1 downto 0);
        CPSEL_FN        : in     vl_logic_vector(2 downto 0);
        KVSEL           : in     vl_logic_vector(1 downto 0);
        FLDD            : in     vl_logic_vector(1 downto 0);
        FORCE_LOCK      : in     vl_logic;
        ATEST_EN        : in     vl_logic;
        DTEST_EN        : in     vl_logic;
        ATEST_SEL       : in     vl_logic;
        DTEST_SEL       : in     vl_logic;
        BP_DVDD12       : in     vl_logic;
        DIVFB           : in     vl_logic;
        CKSEL           : in     vl_logic;
        CK_SWITCH_EN    : in     vl_logic;
        LKD_TOL         : in     vl_logic;
        LKD_HOLD        : in     vl_logic;
        SSEN            : in     vl_logic;
        SSRG            : in     vl_logic_vector(1 downto 0);
        SSDIVH          : in     vl_logic_vector(1 downto 0);
        SSDIVL          : in     vl_logic_vector(7 downto 0);
        BK              : in     vl_logic_vector(1 downto 0);
        CKBAD0          : out    vl_logic;
        CKBAD1          : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of MAX_INPUT_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MIN_INPUT_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MAX_PFD_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MIN_PFD_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MAX_VCO_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MIN_VCO_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MAX_OUTPUT_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of MIN_OUTPUT_PERIOD : constant is 1;
    attribute mti_svvh_generic_type of LOCK_TIME : constant is 1;
end PLL_SIM;
