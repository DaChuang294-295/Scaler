(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/divider_v2.v:3",
  agate_format    = "VLOG"
*)
module mdivider_1(reset, ratio, remainder, error, divisor, dividend);
input reset;
output error;
input  [16:0] divisor;
input  [16:0] dividend;
output [16:0] ratio;
output [16:0] remainder;
reg [16:0] divisor_a;
reg [33:0] shift_dividend;
reg N5;
wire __dbP54, __dbP170, N6, N7, __dbP171, N8, N9, __dbP172, N10, N11, __dbP173,
     N12, N13, __dbP174, N14, N15, __dbP175, N16, N17, __dbP176, N18, N19,
     __dbP177, N20, N21, __dbP178, N22, N23, __dbP179, N24, N25, __dbP180, N26,
     N27, __dbP181, N28, N29, __dbP182, N30, N31, __dbP183, N32, N33, __dbP184,
     N34, N35, __dbP185, N36, n21, n90, n125, n277, n278, n279, n280, n281,
     n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
     n294, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
     n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
     n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
     n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
     n425, n426, n427, n479, n480, n481, n482, n483, n484, n485, n486, n487,
     n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
     n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
     n524, n525, n526, n527, n528, n580, n581, n582, n583, n584, n585, n586,
     n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
     n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
     n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
     n623, n624, n625, n626, n627, n628, n629, n681, n682, n683, n684, n685,
     n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
     n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
     n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
     n722, n723, n724, n725, n726, n727, n728, n729, n730, n782, n783, n784,
     n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
     n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
     n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
     n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n883,
     n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
     n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
     n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
     n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
     n932, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
     n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
     n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
     n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
     n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1085, n1086,
     n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
     n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
     n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
     n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
     n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1186, n1187,
     n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
     n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
     n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
     n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
     n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1287, n1288,
     n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
     n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
     n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
     n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
     n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1388, n1389,
     n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
     n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
     n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
     n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
     n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1489, n1490,
     n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
     n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
     n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
     n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
     n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1590, n1591,
     n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
     n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
     n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
     n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
     n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1691, n1692,
     n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
     n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
     n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
     n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
     n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1792, n1793,
     n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
     n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
     n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
     n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
     n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1963, n1964,
     n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
     n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
     n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
     n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
     n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
     n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
     n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
     n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
     n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
     n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
     n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
     n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
     n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
     n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
     n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
     n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
     n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
     n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
     n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
     n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
     n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
     n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
     n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
     n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
     n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
     n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
     n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
     n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
     n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
     n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
     n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
     n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
     n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
     n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
     n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
     n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
     n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
     n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
     n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
     n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
     n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
     n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
     n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
     n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
     n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
     n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
     n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
     n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
     n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
     n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
     n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
     n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
     n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
     n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
     n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
     n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2541,
     n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
     n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
     n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
     n2572, n2573, n2574, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
     n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
     n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
     n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2883, n2884, n2885,
     n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
     n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
     n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
     n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
     n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/divider_v2.v:3",
  agate_format    = "VLOG"
*)
module mdivider_2(reset, ratio, remainder, error, divisor, dividend);
input reset;
output error;
input  [16:0] divisor;
input  [16:0] dividend;
output [16:0] ratio;
output [16:0] remainder;
reg [16:0] divisor_a;
reg [33:0] shift_dividend;
reg N5;
wire __dbP54, __dbP170, N6, N7, __dbP171, N8, N9, __dbP172, N10, N11, __dbP173,
     N12, N13, __dbP174, N14, N15, __dbP175, N16, N17, __dbP176, N18, N19,
     __dbP177, N20, N21, __dbP178, N22, N23, __dbP179, N24, N25, __dbP180, N26,
     N27, __dbP181, N28, N29, __dbP182, N30, N31, __dbP183, N32, N33, __dbP184,
     N34, N35, __dbP185, N36, n21, n90, n125, n277, n278, n279, n280, n281,
     n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
     n294, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
     n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
     n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
     n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
     n425, n426, n427, n479, n480, n481, n482, n483, n484, n485, n486, n487,
     n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
     n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
     n524, n525, n526, n527, n528, n580, n581, n582, n583, n584, n585, n586,
     n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
     n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
     n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
     n623, n624, n625, n626, n627, n628, n629, n681, n682, n683, n684, n685,
     n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
     n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
     n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
     n722, n723, n724, n725, n726, n727, n728, n729, n730, n782, n783, n784,
     n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
     n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
     n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
     n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n883,
     n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
     n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
     n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
     n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
     n932, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
     n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
     n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
     n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
     n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1085, n1086,
     n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
     n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
     n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
     n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
     n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1186, n1187,
     n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
     n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
     n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
     n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
     n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1287, n1288,
     n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
     n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
     n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
     n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
     n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1388, n1389,
     n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
     n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
     n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
     n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
     n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1489, n1490,
     n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
     n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
     n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
     n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
     n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1590, n1591,
     n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
     n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
     n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
     n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
     n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1691, n1692,
     n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
     n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
     n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
     n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
     n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1792, n1793,
     n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
     n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
     n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
     n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
     n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1963, n1964,
     n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
     n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
     n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
     n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
     n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
     n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
     n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
     n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
     n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
     n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
     n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
     n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
     n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
     n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
     n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
     n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
     n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
     n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
     n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
     n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
     n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
     n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
     n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
     n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
     n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
     n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
     n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
     n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
     n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
     n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
     n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
     n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
     n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
     n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
     n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
     n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
     n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
     n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
     n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
     n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
     n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
     n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
     n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
     n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
     n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
     n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
     n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
     n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
     n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
     n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
     n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
     n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
     n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
     n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
     n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
     n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2541,
     n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
     n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
     n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
     n2572, n2573, n2574, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
     n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
     n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
     n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2883, n2884, n2885,
     n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
     n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
     n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
     n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
     n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/coefcal_v3.v:10",
  agate_format    = "VLOG"
*)
module coefCal_INPUT_RES_WIDTH11_OUTPUT_RES_WIDTH11_SCALE_BITS8(clk, rst, en,
     xBgn, xEnd, yBgn, yEnd, inXRes, inYRes, outXRes, outYRes, kX, kY, inEn,
     iVsyn);
input clk, rst, en, iVsyn;
output inEn;
input  [10:0] xBgn;
input  [10:0] xEnd;
input  [10:0] yBgn;
input  [10:0] yEnd;
input  [10:0] inXRes;
input  [10:0] inYRes;
input  [10:0] outXRes;
input  [10:0] outYRes;
output [7:0] kX;
output [7:0] kY;
reg [8:0] frameRate;
reg [32:0] test;
reg [32:0] working;
reg [16:0] xDividend;
reg [16:0] xDivisor;
reg [16:0] yDividend;
reg [16:0] yDivisor;
wire [16:0] preKX;
wire [16:0] preKY;
reg inEn, work;
wire N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, __dbP50, N13, N15, N16, N17,
     n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
     n19, n20, n21, n22, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
     n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
     n62, n63, n64, n65, n66, n67, n68, n101, n104, n247, n248, n249, n250,
     n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
     n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
     n275, n276, n277, n278, n311, n312, n313, n314, n315, n316, n317, n318,
     n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
     n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
     n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
     n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
     n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
     n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
     n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
     n447, n448, n449, n450, n535, n536, n537, n538, n539, n540, n541, n542,
     n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
     n555, n556, n557, n558, n599, n600, n601, n602, n603, n604, n605, n606,
     n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
     n619, n620, n621, n622, n625, n626, n627, n628, n629, n916, n917, n918,
     n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
     n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
     n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
     n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
     n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
     n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
     n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
     n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
     n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
     n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
     n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
     n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
     n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
     n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
     n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
     n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
     n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
     n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
     n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
     n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
     n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
     n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
     n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
     n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
     n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
     n1183, n1184, n1185, n1186, n1187, n1188;
    mdivider_1 divide_inst1 (.reset(rst), .ratio({preKX[16:0]}), .divisor({xDivisor[16:0]}),
        .dividend({xDividend[16:0]}));
    mdivider_2 divide_inst2 (.reset(rst), .ratio({preKY[16:0]}), .divisor({yDivisor[16:0]}),
        .dividend({yDividend[16:0]}));

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/inputCtrl.v:9",
  agate_format    = "VLOG"
*)
module inputCtrl_DATA_WIDTH16_INPUT_RES_WIDTH11_SCALE_FRAC_WIDTH6_SCALE_INT_WIDTH2_ADDRESS_WIDTH11(clk,
     rst, xBgn, xEnd, yBgn, yEnd, dInEn, dIn, iHsyn, iVsyn, En, kX, kY,
     ramWrtAddr, ramWrtEn, dataOut, jmp);
input clk, rst, dInEn, iHsyn, iVsyn, En;
output ramWrtEn, jmp;
input  [10:0] xBgn;
input  [10:0] xEnd;
input  [10:0] yBgn;
input  [10:0] yEnd;
input  [15:0] dIn;
input  [7:0] kX;
input  [7:0] kY;
output [10:0] ramWrtAddr;
output [15:0] dataOut;
reg [15:0] dataOut;
reg [10:0] ramWrtAddr;
reg [10:0] xAddress;
reg [16:0] xCal;
reg [10:0] yAddress;
reg [16:0] yCal;
wire [7:0] xAdder;
wire [10:0] xNxtAddress;
wire [16:0] xNxtCal;
wire [7:0] yAdder;
wire [10:0] yNxtAddress;
wire [16:0] yNxtCal;
reg jmp, ramWrtEn, xPreEn, yPreEn;
wire boundEn, trueEn, xBgnEn, xEn, xEndEn, xRst, xThisEn, yBgnEn, yEn, yEndEn,
     yRst, yThisEn, __dbP19, __dbP36, N1, N2, N3, N4, __dbP109, __dbP174,
     __dbP239, __dbP304, N5, n19, n20, n45, n46, n140, n141, n142, n143, n144,
     n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
     n157, n158, n159, n160, n204, n205, n206, n207, n208, n209, n210, n211,
     n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
     n224, n225, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
     n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
     n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n388, n389,
     n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
     n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
     n414, n415, n416, n417, n418, n419, n485, n486, n487, n488, n489, n490,
     n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
     n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
     n515, n516, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
     n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
     n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n679, n680,
     n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
     n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
     n705, n706, n707, n708, n709, n710, n776, n777, n778, n779, n780, n781,
     n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
     n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
     n806, n845, n928, n972, n973, n974, n975, n976, n977, n978, n979, n980,
     n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
     n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
     n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
     n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
     n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
     n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
     n1073, n1074, n1075, n1076, n1077, n1078, n1137, n1138, n1139, n1140,
     n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
     n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
     n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
     n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
     n1181, n1182, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
     n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
     n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
     n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
     n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
     n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
     n1299, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
     n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
     n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
     n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
     n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
     n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
     n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
     n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
     n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662;

endmodule

(*
  agate_file_name = "/cygdrive/F/capital_micro/primace7.3/ast_frontend//../data/lib/syn_black_box_m7s.v:427",
  agate_format    = "VLOG"
*)
module M7S_EMB18K(wfull, wfull_almost, rempty, rempty_almost, overflow, wr_ack,
     underflow, rd_ack, rd_ha, rd_la, c1r4_q, c1r3_q, c1r2_q, c1r1_q, c1r4_aa,
     c1r4_ab, c1r4_cea, c1r4_ceb, c1r4_clka, c1r4_clkb, c1r4_da, c1r4_db,
     c1r4_rstna, c1r4_rstnb, c1r4_wea, c1r4_web, c1r3_aa, c1r3_ab, c1r3_cea,
     c1r3_ceb, c1r3_clka, c1r3_clkb, c1r3_da, c1r3_db, c1r3_rstna, c1r3_rstnb,
     c1r3_wea, c1r3_web, c1r2_aa, c1r2_ab, c1r2_cea, c1r2_ceb, c1r2_clka,
     c1r2_clkb, c1r2_da, c1r2_db, c1r2_rstna, c1r2_rstnb, c1r2_wea, c1r2_web,
     c1r1_aa, c1r1_ab, c1r1_cea, c1r1_ceb, c1r1_clka, c1r1_clkb, c1r1_da,
     c1r1_db, c1r1_rstna, c1r1_rstnb, c1r1_wea, c1r1_web, cea, ceb, fifo_clr,
     wr_req_n, rd_req_n, haa, hab, wea, web);
input c1r4_cea, c1r4_ceb, c1r4_clka, c1r4_clkb, c1r4_rstna, c1r4_rstnb,
     c1r4_wea, c1r4_web, c1r3_cea, c1r3_ceb, c1r3_clka, c1r3_clkb, c1r3_rstna,
     c1r3_rstnb, c1r3_wea, c1r3_web, c1r2_cea, c1r2_ceb, c1r2_clka, c1r2_clkb,
     c1r2_rstna, c1r2_rstnb, c1r2_wea, c1r2_web, c1r1_cea, c1r1_ceb, c1r1_clka,
     c1r1_clkb, c1r1_rstna, c1r1_rstnb, c1r1_wea, c1r1_web, cea, ceb, fifo_clr,
     wr_req_n, rd_req_n, wea, web;
output wfull, wfull_almost, rempty, rempty_almost, overflow, wr_ack, underflow,
     rd_ack;
input  [11:0] c1r4_aa;
input  [11:0] c1r4_ab;
input  [17:0] c1r4_da;
input  [17:0] c1r4_db;
input  [11:0] c1r3_aa;
input  [11:0] c1r3_ab;
input  [17:0] c1r3_da;
input  [17:0] c1r3_db;
input  [11:0] c1r2_aa;
input  [11:0] c1r2_ab;
input  [17:0] c1r2_da;
input  [17:0] c1r2_db;
input  [11:0] c1r1_aa;
input  [11:0] c1r1_ab;
input  [17:0] c1r1_da;
input  [17:0] c1r1_db;
input  [1:0] haa;
input  [1:0] hab;
output [1:0] rd_ha;
output [5:0] rd_la;
output [17:0] c1r4_q;
output [17:0] c1r3_q;
output [17:0] c1r2_q;
output [17:0] c1r1_q;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/emb_16_2k.v:14",
  agate_format    = "VLOG"
*)
module emb_16_2k_1(clka, cea, wea, aa, da, qa, clkb, ceb, web, ab, db, qb);
input clka, cea, wea, clkb, ceb, web;
input  [10:0] aa;
input  [15:0] da;
input  [10:0] ab;
input  [15:0] db;
output [15:0] qa;
output [15:0] qb;
reg [0:0] aa_reg;
reg [0:0] ab_reg;
wire [8:0] qa0;
wire [8:0] qa1;
wire [8:0] qa2;
wire [8:0] qa3;
wire [8:0] qa4;
wire [8:0] qa5;
wire [8:0] qa6;
wire [8:0] qa7;
wire [8:0] qb0;
wire [8:0] qb1;
wire [8:0] qb2;
wire [8:0] qb3;
wire [8:0] qb4;
wire [8:0] qb5;
wire [8:0] qb6;
wire [8:0] qb7;
wire n3, n52, n102, n105, n113, n114, n115, n116, n117, n118, n119, n120, n121,
     n122, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
     n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
     n152, n153, n154, n159, n160, n161, n162, n163, n164, n165, n166, n167,
     n168, n169, n170, n171, n172, n173, n174, n199, n200, n201, n202, n203,
     n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n219,
     n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
     n232, n233, n234, n259, n260, n261, n262, n263, n264, n265, n266, n267,
     n268, n269, n270, n271, n272, n273, n274, n279, n280, n281, n282, n283,
     n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n319,
     n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
     n332, n333, n334, n339, n340, n341, n342, n343, n344, n345, n346, n347,
     n348, n349, n350, n351, n352, n353, n354, n376, n379, n387, n388, n389,
     n390, n391, n392, n393, n394, n395, n396, n401, n402, n403, n404, n405,
     n406, n407, n408, n409, n410, n413, n414, n415, n416, n417, n418, n419,
     n420, n421, n422, n423, n424, n425, n426, n427, n428, n433, n434, n435,
     n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
     n448, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
     n484, n485, n486, n487, n488, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n533, n534, n535,
     n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
     n548, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
     n564, n565, n566, n567, n568, n593, n594, n595, n596, n597, n598, n599,
     n600, n601, n602, n603, n604, n605, n606, n607, n608, n613, n614, n615,
     n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
     n628, n649, n650, n889, n890;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/emb_16_2k.v:14",
  agate_format    = "VLOG"
*)
module emb_16_2k_2(clka, cea, wea, aa, da, qa, clkb, ceb, web, ab, db, qb);
input clka, cea, wea, clkb, ceb, web;
input  [10:0] aa;
input  [15:0] da;
input  [10:0] ab;
input  [15:0] db;
output [15:0] qa;
output [15:0] qb;
reg [0:0] aa_reg;
reg [0:0] ab_reg;
wire [8:0] qa0;
wire [8:0] qa1;
wire [8:0] qa2;
wire [8:0] qa3;
wire [8:0] qa4;
wire [8:0] qa5;
wire [8:0] qa6;
wire [8:0] qa7;
wire [8:0] qb0;
wire [8:0] qb1;
wire [8:0] qb2;
wire [8:0] qb3;
wire [8:0] qb4;
wire [8:0] qb5;
wire [8:0] qb6;
wire [8:0] qb7;
wire n3, n52, n102, n105, n113, n114, n115, n116, n117, n118, n119, n120, n121,
     n122, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
     n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
     n152, n153, n154, n159, n160, n161, n162, n163, n164, n165, n166, n167,
     n168, n169, n170, n171, n172, n173, n174, n199, n200, n201, n202, n203,
     n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n219,
     n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
     n232, n233, n234, n259, n260, n261, n262, n263, n264, n265, n266, n267,
     n268, n269, n270, n271, n272, n273, n274, n279, n280, n281, n282, n283,
     n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n319,
     n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
     n332, n333, n334, n339, n340, n341, n342, n343, n344, n345, n346, n347,
     n348, n349, n350, n351, n352, n353, n354, n376, n379, n387, n388, n389,
     n390, n391, n392, n393, n394, n395, n396, n401, n402, n403, n404, n405,
     n406, n407, n408, n409, n410, n413, n414, n415, n416, n417, n418, n419,
     n420, n421, n422, n423, n424, n425, n426, n427, n428, n433, n434, n435,
     n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
     n448, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
     n484, n485, n486, n487, n488, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n533, n534, n535,
     n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
     n548, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
     n564, n565, n566, n567, n568, n593, n594, n595, n596, n597, n598, n599,
     n600, n601, n602, n603, n604, n605, n606, n607, n608, n613, n614, n615,
     n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
     n628, n649, n650, n889, n890;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/emb_16_2k.v:14",
  agate_format    = "VLOG"
*)
module emb_16_2k_3(clka, cea, wea, aa, da, qa, clkb, ceb, web, ab, db, qb);
input clka, cea, wea, clkb, ceb, web;
input  [10:0] aa;
input  [15:0] da;
input  [10:0] ab;
input  [15:0] db;
output [15:0] qa;
output [15:0] qb;
reg [0:0] aa_reg;
reg [0:0] ab_reg;
wire [8:0] qa0;
wire [8:0] qa1;
wire [8:0] qa2;
wire [8:0] qa3;
wire [8:0] qa4;
wire [8:0] qa5;
wire [8:0] qa6;
wire [8:0] qa7;
wire [8:0] qb0;
wire [8:0] qb1;
wire [8:0] qb2;
wire [8:0] qb3;
wire [8:0] qb4;
wire [8:0] qb5;
wire [8:0] qb6;
wire [8:0] qb7;
wire n3, n52, n102, n105, n113, n114, n115, n116, n117, n118, n119, n120, n121,
     n122, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
     n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
     n152, n153, n154, n159, n160, n161, n162, n163, n164, n165, n166, n167,
     n168, n169, n170, n171, n172, n173, n174, n199, n200, n201, n202, n203,
     n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n219,
     n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
     n232, n233, n234, n259, n260, n261, n262, n263, n264, n265, n266, n267,
     n268, n269, n270, n271, n272, n273, n274, n279, n280, n281, n282, n283,
     n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n319,
     n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
     n332, n333, n334, n339, n340, n341, n342, n343, n344, n345, n346, n347,
     n348, n349, n350, n351, n352, n353, n354, n376, n379, n387, n388, n389,
     n390, n391, n392, n393, n394, n395, n396, n401, n402, n403, n404, n405,
     n406, n407, n408, n409, n410, n413, n414, n415, n416, n417, n418, n419,
     n420, n421, n422, n423, n424, n425, n426, n427, n428, n433, n434, n435,
     n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
     n448, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
     n484, n485, n486, n487, n488, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n533, n534, n535,
     n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
     n548, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
     n564, n565, n566, n567, n568, n593, n594, n595, n596, n597, n598, n599,
     n600, n601, n602, n603, n604, n605, n606, n607, n608, n613, n614, n615,
     n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
     n628, n649, n650, n889, n890;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/emb_16_2k.v:14",
  agate_format    = "VLOG"
*)
module emb_16_2k_4(clka, cea, wea, aa, da, qa, clkb, ceb, web, ab, db, qb);
input clka, cea, wea, clkb, ceb, web;
input  [10:0] aa;
input  [15:0] da;
input  [10:0] ab;
input  [15:0] db;
output [15:0] qa;
output [15:0] qb;
reg [0:0] aa_reg;
reg [0:0] ab_reg;
wire [8:0] qa0;
wire [8:0] qa1;
wire [8:0] qa2;
wire [8:0] qa3;
wire [8:0] qa4;
wire [8:0] qa5;
wire [8:0] qa6;
wire [8:0] qa7;
wire [8:0] qb0;
wire [8:0] qb1;
wire [8:0] qb2;
wire [8:0] qb3;
wire [8:0] qb4;
wire [8:0] qb5;
wire [8:0] qb6;
wire [8:0] qb7;
wire n3, n52, n102, n105, n113, n114, n115, n116, n117, n118, n119, n120, n121,
     n122, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n139,
     n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
     n152, n153, n154, n159, n160, n161, n162, n163, n164, n165, n166, n167,
     n168, n169, n170, n171, n172, n173, n174, n199, n200, n201, n202, n203,
     n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n219,
     n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
     n232, n233, n234, n259, n260, n261, n262, n263, n264, n265, n266, n267,
     n268, n269, n270, n271, n272, n273, n274, n279, n280, n281, n282, n283,
     n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n319,
     n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
     n332, n333, n334, n339, n340, n341, n342, n343, n344, n345, n346, n347,
     n348, n349, n350, n351, n352, n353, n354, n376, n379, n387, n388, n389,
     n390, n391, n392, n393, n394, n395, n396, n401, n402, n403, n404, n405,
     n406, n407, n408, n409, n410, n413, n414, n415, n416, n417, n418, n419,
     n420, n421, n422, n423, n424, n425, n426, n427, n428, n433, n434, n435,
     n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
     n448, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
     n484, n485, n486, n487, n488, n493, n494, n495, n496, n497, n498, n499,
     n500, n501, n502, n503, n504, n505, n506, n507, n508, n533, n534, n535,
     n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
     n548, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
     n564, n565, n566, n567, n568, n593, n594, n595, n596, n597, n598, n599,
     n600, n601, n602, n603, n604, n605, n606, n607, n608, n613, n614, n615,
     n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
     n628, n649, n650, n889, n890;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/ramFifo.v:9",
  agate_format    = "VLOG"
*)
module ramFifo_DATA_WIDTH16_ADDRESS_WIDTH11(clka, clkb, rst, advanceRead1,
     advanceRead2, advanceWrite, writeData, writeAddress, writeEnable,
     fillCount, readData00, readData01, readData10, readData11, readAddress00,
     readAddress01, readAddress10, readAddress11);
input clka, clkb, rst, advanceRead1, advanceRead2, advanceWrite, writeEnable;
input  [15:0] writeData;
input  [10:0] writeAddress;
input  [10:0] readAddress00;
input  [10:0] readAddress01;
input  [10:0] readAddress10;
input  [10:0] readAddress11;
output [2:0] fillCount;
output [15:0] readData00;
output [15:0] readData01;
output [15:0] readData10;
output [15:0] readData11;
wire [15:0] \ramDataOutA[0] ;
wire [15:0] \ramDataOutA[10] ;
wire [15:0] \ramDataOutA[11] ;
wire [15:0] \ramDataOutA[12] ;
wire [15:0] \ramDataOutA[13] ;
wire [15:0] \ramDataOutA[14] ;
wire [15:0] \ramDataOutA[15] ;
wire [15:0] \ramDataOutA[1] ;
wire [15:0] \ramDataOutA[2] ;
wire [15:0] \ramDataOutA[3] ;
wire [15:0] \ramDataOutA[4] ;
wire [15:0] \ramDataOutA[5] ;
wire [15:0] \ramDataOutA[6] ;
wire [15:0] \ramDataOutA[7] ;
wire [15:0] \ramDataOutA[8] ;
wire [15:0] \ramDataOutA[9] ;
wire [15:0] \ramDataOutB[0] ;
wire [15:0] \ramDataOutB[10] ;
wire [15:0] \ramDataOutB[11] ;
wire [15:0] \ramDataOutB[12] ;
wire [15:0] \ramDataOutB[13] ;
wire [15:0] \ramDataOutB[14] ;
wire [15:0] \ramDataOutB[15] ;
wire [15:0] \ramDataOutB[1] ;
wire [15:0] \ramDataOutB[2] ;
wire [15:0] \ramDataOutB[3] ;
wire [15:0] \ramDataOutB[4] ;
wire [15:0] \ramDataOutB[5] ;
wire [15:0] \ramDataOutB[6] ;
wire [15:0] \ramDataOutB[7] ;
wire [15:0] \ramDataOutB[8] ;
wire [15:0] \ramDataOutB[9] ;
wire [10:0] readAddressA0;
wire [10:0] readAddressA1;
wire [10:0] readAddressB0;
wire [10:0] readAddressB1;
wire [10:0] readAddressC0;
wire [10:0] readAddressC1;
wire [10:0] readAddressD0;
wire [10:0] readAddressD1;
wire [3:0] readSelect;
wire [3:0] readSelect0;
wire [3:0] readSelect1;
wire [3:0] writeSelect;
wire clka0, clka1, clka2, clka3, N5, N6, N7, N8, n159, n160, n161, n162, n163,
     n164, n165, n166, n167, n168, n169, n171, n269, n270, n271, n272, n273,
     n274, n275, n276, n277, n278, n279, n281, n379, n380, n381, n382, n383,
     n384, n385, n386, n387, n388, n389, n391, n489, n490, n491, n492, n493,
     n494, n495, n496, n497, n498, n499, n501, n667, n668, n669, n670, n671,
     n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
     n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
     n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
     n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
     n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
     n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
     n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
     n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
     n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
     n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
     n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
     n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
     n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
     n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
     n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
     n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
     n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
     n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
     n888, n889, n890, n907, n908, n909, n910, n911, n912, n913, n914, n915,
     n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
     n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
     n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
     n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
     n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
     n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
     n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
     n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
     n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
     n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
     n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
     n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
     n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
     n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
     n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
     n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
     n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
     n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
     n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
     n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
     n1130, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
     n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
     n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
     n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
     n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
     n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
     n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
     n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
     n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
     n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
     n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
     n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
     n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
     n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
     n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
     n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
     n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
     n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
     n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
     n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
     n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
     n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
     n1366, n1367, n1368, n1369, n1370, n1387, n1388, n1389, n1390, n1391,
     n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
     n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
     n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
     n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
     n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
     n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
     n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
     n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
     n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
     n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
     n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
     n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
     n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
     n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
     n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
     n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
     n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
     n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
     n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
     n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
     n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
     n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1691,
     n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
     n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
     n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
     n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
     n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
     n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
     n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
     n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
     n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
     n1782, n1783, n1784, n1785, n1786, n1819, n1820, n1821, n1822, n1823,
     n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
     n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
     n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1869, n1870, n1871,
     n1872, n1873, n1874, n1875, n1876, n1890, n1891, n1892, n1893, n1928,
     n1929, n1930, n1931, n1932, n1933, n1951, n1952, n1953, n1954, n1955,
     n1956, n1957, n1958, n1959;
    emb_16_2k_1 ram_inst_0 (.clka(clka0), .cea(), .wea(n171), .aa({n169,
        n168, n167, n166, n165, n164, n163, n162, n161, n160, n159}), .da({writeData[15:0]}),
        .qa({\ramDataOutA[1] [15:0]}), .clkb(clkb), .ceb(), .web(),
        .ab({readAddressA1[10:0]}), .db({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .qb({\ramDataOutB[1] [15:0]}));
    emb_16_2k_2 ram_inst_1 (.clka(clka1), .cea(), .wea(n281), .aa({n279,
        n278, n277, n276, n275, n274, n273, n272, n271, n270, n269}), .da({writeData[15:0]}),
        .qa({\ramDataOutA[2] [15:0]}), .clkb(clkb), .ceb(), .web(),
        .ab({readAddressB1[10:0]}), .db({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .qb({\ramDataOutB[2] [15:0]}));
    emb_16_2k_3 ram_inst_2 (.clka(clka2), .cea(), .wea(n391), .aa({n389,
        n388, n387, n386, n385, n384, n383, n382, n381, n380, n379}), .da({writeData[15:0]}),
        .qa({\ramDataOutA[4] [15:0]}), .clkb(clkb), .ceb(), .web(),
        .ab({readAddressC1[10:0]}), .db({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .qb({\ramDataOutB[4] [15:0]}));
    emb_16_2k_4 ram_inst_3 (.clka(clka3), .cea(), .wea(n501), .aa({n499,
        n498, n497, n496, n495, n494, n493, n492, n491, n490, n489}), .da({writeData[15:0]}),
        .qa({\ramDataOutA[8] [15:0]}), .clkb(clkb), .ceb(), .web(),
        .ab({readAddressD1[10:0]}), .db({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .qb({\ramDataOutB[8] [15:0]}));

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/Cal_v1.v:11",
  agate_format    = "VLOG"
*)
module Cal_DATA_WIDTH16_ADDRESS_WIDTH11_SCALE_FRAC_WIDTH6_SCALE_INT_WIDTH2_INPUT_RES_WIDTH11_OUTPUT_RES_WIDTH11(clk,
     rst, ramAddrIn, ramData00, ramData01, ramData10, ramData11, fifoNum, kX,
     kY, inXNum, inYNum, outXRes, outYRes, HS, VS, dOutEn, jmp1, jmp2,
     ramRdAddr00, ramRdAddr01, ramRdAddr10, ramRdAddr11, dOut);
input clk, rst;
output HS, VS, dOutEn, jmp1, jmp2;
input  [10:0] ramAddrIn;
input  [15:0] ramData00;
input  [15:0] ramData01;
input  [15:0] ramData10;
input  [15:0] ramData11;
input  [1:0] fifoNum;
input  [7:0] kX;
input  [7:0] kY;
input  [10:0] inXNum;
input  [10:0] inYNum;
input  [10:0] outXRes;
input  [10:0] outYRes;
output [10:0] ramRdAddr00;
output [10:0] ramRdAddr01;
output [10:0] ramRdAddr10;
output [10:0] ramRdAddr11;
output [15:0] dOut;
reg [10:0] ramRdAddr;
reg [16:0] u;
reg [5:0] uPreF;
reg [16:0] v;
reg [10:0] xAddress;
reg [10:0] yAddress;
wire [6:0] F00;
wire [11:0] F00B00;
wire [12:0] F00G00;
wire [11:0] F00R00;
wire [5:0] F01;
wire [10:0] F01B01;
wire [11:0] F01G01;
wire [10:0] F01R01;
wire [5:0] F10;
wire [10:0] F10B10;
wire [11:0] F10G10;
wire [10:0] F10R10;
wire [5:0] F11;
wire [10:0] F11B11;
wire [11:0] F11G11;
wire [10:0] F11R11;
wire [4:0] dB00;
wire [4:0] dB01;
wire [4:0] dB10;
wire [4:0] dB11;
wire [4:0] dBout;
wire [5:0] dG00;
wire [5:0] dG01;
wire [5:0] dG10;
wire [5:0] dG11;
wire [5:0] dGout;
wire [4:0] dR00;
wire [4:0] dR01;
wire [4:0] dR10;
wire [4:0] dR11;
wire [4:0] dRout;
wire [15:0] data00;
wire [15:0] data01;
wire [15:0] data10;
wire [15:0] data11;
wire [11:0] preuv;
wire [2:0] uDistance;
wire [5:0] uF;
wire [10:0] uI;
wire [2:0] uIK;
wire [16:0] uNxt;
wire [2:0] uNxtIK;
wire [5:0] uv;
wire [2:0] vDistance;
wire [5:0] vF;
wire [10:0] vI;
wire [2:0] vIK;
wire [16:0] vNxt;
wire [2:0] vNxtIK;
wire [1:0] xAddrDistance;
wire [1:0] yAddrDistance;
reg HS, VSNormal, enforceJmp, jmp1Normal, jmp2Normal;
wire enCal, inXBound, inYBound, mode, outXBoundEn, outXLowEn, outXUpEn,
     outYBoundEn, outYLowEn, outYUpEn, workEn, N1, N2, __dbP67, N3, N4,
     __dbP132, __dbP167, __dbP360, __dbP425, __dbP522, __dbP587, __dbP652,
     __dbP717, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
     N19, N20, N21, N22, n55, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99,
     n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
     n112, n113, n114, n115, n116, n117, n118, n119, n172, n177, n210, n276,
     n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
     n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
     n301, n302, n303, n304, n305, n306, n339, n405, n406, n407, n408, n409,
     n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
     n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
     n434, n435, n468, n534, n535, n536, n537, n538, n539, n540, n541, n542,
     n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
     n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n631,
     n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
     n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
     n656, n657, n658, n659, n660, n661, n695, n761, n762, n763, n764, n765,
     n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
     n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
     n790, n791, n792, n858, n859, n860, n861, n862, n863, n864, n865, n866,
     n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
     n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n890, n956,
     n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
     n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
     n981, n982, n983, n984, n985, n986, n987, n1053, n1054, n1055, n1056,
     n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
     n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
     n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
     n1087, n1088, n1089, n1157, n1190, n1223, n1224, n1225, n1226, n1227,
     n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
     n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
     n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1266, n1267, n1268,
     n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
     n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1353,
     n1354, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
     n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
     n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
     n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
     n1426, n1427, n1428, n1429, n1430, n1495, n1497, n1498, n1499, n1500,
     n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
     n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
     n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1536,
     n1537, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
     n1610, n1611, n1612, n1613, n1614, n1773, n1774, n1775, n1776, n1777,
     n1778, n1779, n1780, n1781, n1782, n1788, n1789, n1790, n1791, n1792,
     n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1806, n1807, n1808,
     n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1822, n1826, n1828,
     n1829, n1830, n1877, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
     n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
     n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
     n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
     n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
     n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2040,
     n2041, n2042, n2043, n2044, n2045, n2134, n2135, n2136, n2137, n2138,
     n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
     n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
     n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
     n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
     n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
     n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
     n2199, n2200, n2201, n2202, n2203, n2204, n2237, n2238, n2939, n2940,
     n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
     n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
     n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
     n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
     n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
     n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
     n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
     n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
     n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
     n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
     n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
     n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
     n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
     n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
     n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
     n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
     n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
     n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
     n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
     n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
     n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
     n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
     n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
     n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
     n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
     n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
     n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
     n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
     n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
     n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
     n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
     n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
     n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
     n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
     n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
     n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
     n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
     n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319;

endmodule

(*
  agate_file_name = "/cygdrive/f/capital_micro/primace7.3/bin/dachuang/final_scaler_v3/outputs/../src/scaler1.0.v:8",
  agate_format    = "VLOG"
*)
module scaler(clka, clkb, rst, en, iHsyn, iVsyn, dIn, dInEn, dOut, dOutEn, HS,
     VS, xBgn, xEnd, yBgn, yEnd, inYRes, inXRes, outYRes, outXRes);
input clka, clkb, rst, en, iHsyn, iVsyn, dInEn;
output dOutEn, HS, VS;
input  [15:0] dIn;
input  [10:0] xBgn;
input  [10:0] xEnd;
input  [10:0] yBgn;
input  [10:0] yEnd;
input  [10:0] inYRes;
input  [10:0] inXRes;
input  [11:0] outYRes;
input  [11:0] outXRes;
output [15:0] dOut;
wire [2:0] fifoNum;
wire [7:0] kX;
wire [7:0] kY;
wire [15:0] ramData;
wire [15:0] ramData00;
wire [15:0] ramData01;
wire [15:0] ramData10;
wire [15:0] ramData11;
wire [10:0] ramRdAddr00;
wire [10:0] ramRdAddr01;
wire [10:0] ramRdAddr10;
wire [10:0] ramRdAddr11;
wire [10:0] ramWrtAddr;
wire inEn, jmp, jmp1, jmp2, ramWrtEn, N156, N158, n3, n4, n5, n6, n7, n8, n9,
     n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
     n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n67, n68, n69, n70, n71,
     n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
     n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
     n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
     n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
     n125, n126, n127, n128, n129, n130, n163, n164, n165, n166, n167, n168,
     n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
     n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
     n193, n194;
    coefCal_INPUT_RES_WIDTH11_OUTPUT_RES_WIDTH11_SCALE_BITS8 coefcal1 (.clk(clka),
        .rst(rst), .en(en), .xBgn({xBgn[10:0]}), .xEnd({xEnd[10:0]}), .yBgn({yBgn[10:0]}),
        .yEnd({yEnd[10:0]}), .inXRes({inXRes[10:0]}), .inYRes({inYRes[10:0]}),
        .outXRes({outXRes[10:0]}), .outYRes({outYRes[10:0]}), .kX({kX[7:0]}),
        .kY({kY[7:0]}), .inEn(inEn), .iVsyn(iVsyn));
    defparam coefcal1.INPUT_RES_WIDTH = 11;
    defparam coefcal1.OUTPUT_RES_WIDTH = 11;
    defparam coefcal1.SCALE_BITS = 8;
    inputCtrl_DATA_WIDTH16_INPUT_RES_WIDTH11_SCALE_FRAC_WIDTH6_SCALE_INT_WIDTH2_ADDRESS_WIDTH11 inputctrl1 (.clk(clka),
        .rst(rst), .xBgn({xBgn[10:0]}), .xEnd({xEnd[10:0]}), .yBgn({yBgn[10:0]}),
        .yEnd({yEnd[10:0]}), .dInEn(dInEn), .dIn({dIn[15:0]}), .iHsyn(iHsyn),
        .iVsyn(iVsyn), .En(inEn), .kX({kX[7:0]}), .kY({kY[7:0]}), .ramWrtAddr({ramWrtAddr[10:0]}),
        .ramWrtEn(ramWrtEn), .dataOut({ramData[15:0]}), .jmp(jmp));
    defparam inputctrl1.DATA_WIDTH = 16;
    defparam inputctrl1.INPUT_RES_WIDTH = 11;
    defparam inputctrl1.SCALE_FRAC_WIDTH = 6;
    defparam inputctrl1.SCALE_INT_WIDTH = 2;
    defparam inputctrl1.ADDRESS_WIDTH = 11;
    ramFifo_DATA_WIDTH16_ADDRESS_WIDTH11 fifo1 (.clka(clka), .clkb(clkb),
        .rst(rst), .advanceRead1(jmp1), .advanceRead2(jmp2), .advanceWrite(jmp),
        .writeData({ramData[15:0]}), .writeAddress({ramWrtAddr[10:0]}), .writeEnable(ramWrtEn),
        .fillCount({fifoNum[2:0]}), .readData00({ramData00[15:0]}), .readData01({ramData01[15:0]}),
        .readData10({ramData10[15:0]}), .readData11({ramData11[15:0]}), .readAddress00({ramRdAddr00[10:0]}),
        .readAddress01({ramRdAddr01[10:0]}), .readAddress10({ramRdAddr10[10:0]}),
        .readAddress11({ramRdAddr11[10:0]}));
    defparam fifo1.DATA_WIDTH = 16;
    defparam fifo1.ADDRESS_WIDTH = 11;
    Cal_DATA_WIDTH16_ADDRESS_WIDTH11_SCALE_FRAC_WIDTH6_SCALE_INT_WIDTH2_INPUT_RES_WIDTH11_OUTPUT_RES_WIDTH11 cal1 (.clk(clkb),
        .rst(rst), .ramAddrIn({ramData[10:0]}), .ramData00({ramData00[15:0]}),
        .ramData01({ramData01[15:0]}), .ramData10({ramData10[15:0]}), .ramData11({ramData11[15:0]}),
        .fifoNum({fifoNum[1:0]}), .kX({kX[7:0]}), .kY({kY[7:0]}), .inXNum({n77,
        n76, n75, n74, n73, n72, n71, n70, n69, n68, n67}), .inYNum({n173,
        n172, n171, n170, n169, n168, n167, n166, n165, n164, n163}), .outXRes({outXRes[10:0]}),
        .outYRes({outYRes[10:0]}), .HS(HS), .VS(VS), .dOutEn(dOutEn), .jmp1(jmp1),
        .jmp2(jmp2), .ramRdAddr00({ramRdAddr00[10:0]}), .ramRdAddr01({ramRdAddr01[10:0]}),
        .ramRdAddr10({ramRdAddr10[10:0]}), .ramRdAddr11({ramRdAddr11[10:0]}),
        .dOut({dOut[15:0]}));
    defparam cal1.DATA_WIDTH = 16;
    defparam cal1.ADDRESS_WIDTH = 11;
    defparam cal1.SCALE_INT_WIDTH = 2;
    defparam cal1.SCALE_FRAC_WIDTH = 6;
    defparam cal1.INPUT_RES_WIDTH = 11;
    defparam cal1.OUTPUT_RES_WIDTH = 11;

endmodule

