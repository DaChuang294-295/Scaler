library verilog;
use verilog.vl_types.all;
entity M7A_IO_DDRSG is
    generic(
        cfg_nc          : vl_logic := Hi0;
        cfg_use_cal1    : vl_logic := Hi0;
        odt_cfg         : vl_logic := Hi0;
        ns_lv_cfg       : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pdr_cfg         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ndr_cfg         : vl_logic_vector(0 to 4) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        keep_cfg        : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        term_pu_en      : vl_logic := Hi0;
        term_pd_en      : vl_logic := Hi0;
        rx_dig_en_cfg   : vl_logic := Hi0;
        rx_hstl_sstl_en_cfg: vl_logic := Hi0;
        tpd_cfg         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        tpu_cfg         : vl_logic_vector(0 to 7) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        cfg_trm         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        cfg_trm_sel     : vl_logic := Hi0;
        in_del          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        out_del         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        cfg_test_en     : vl_logic := Hi0;
        cfg_userio_en   : vl_logic := Hi0;
        cfg_use_cal0    : vl_logic := Hi0;
        cfg_fclk_inv    : vl_logic := Hi0;
        cfg_gsclk_inv   : vl_logic := Hi0;
        cfg_gsclk90_inv : vl_logic := Hi0;
        cfg_gsclk180_inv: vl_logic := Hi0;
        cfg_gsclk270_inv: vl_logic := Hi0;
        cfg_fclk_gate_sel: vl_logic := Hi0;
        cfg_sclk_gate_sel: vl_logic := Hi0;
        cfg_sclk_en     : vl_logic := Hi0;
        cfg_fclk_en     : vl_logic := Hi0;
        cfg_rstn_inv    : vl_logic := Hi0;
        cfg_oen_rstn_en : vl_logic := Hi0;
        cfg_od_rstn_en  : vl_logic := Hi0;
        cfg_id_rstn_en  : vl_logic := Hi0;
        cfg_setn_inv    : vl_logic := Hi0;
        cfg_oen_setn_en : vl_logic := Hi0;
        cfg_od_setn_en  : vl_logic := Hi0;
        cfg_id_setn_en  : vl_logic := Hi0;
        cfg_ddr         : vl_logic := Hi0;
        cfg_id_sel      : vl_logic := Hi0;
        cfg_oen_inv     : vl_logic := Hi0;
        cfg_oen_sel     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_dqs         : vl_logic := Hi0;
        cfg_txd0_inv    : vl_logic := Hi0;
        cfg_txd1_inv    : vl_logic := Hi0;
        cfg_d_en        : vl_logic := Hi0;
        cfg_clkout_sel  : vl_logic := Hi0;
        cfg_sclk_out    : vl_logic := Hi0;
        cfg_od_sel      : vl_logic_vector(0 to 1) := (Hi0, Hi0)
    );
    port(
        id_q            : out    vl_logic_vector(1 downto 0);
        NDR_in          : in     vl_logic_vector(4 downto 0);
        PDR_in          : in     vl_logic_vector(4 downto 0);
        TPD_in          : in     vl_logic_vector(7 downto 0);
        TPU_in          : in     vl_logic_vector(7 downto 0);
        clk_en          : in     vl_logic;
        clkpol          : in     vl_logic;
        dqsr90          : in     vl_logic;
        gsclk270_in     : in     vl_logic;
        gsclk180_in     : in     vl_logic;
        gsclk90_in      : in     vl_logic;
        gsclk_in        : in     vl_logic;
        od_d            : in     vl_logic_vector(1 downto 0);
        oen             : in     vl_logic;
        clk             : in     vl_logic;
        rstn            : in     vl_logic;
        setn            : in     vl_logic;
        PAD             : inout  vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of cfg_nc : constant is 1;
    attribute mti_svvh_generic_type of cfg_use_cal1 : constant is 1;
    attribute mti_svvh_generic_type of odt_cfg : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_cfg : constant is 1;
    attribute mti_svvh_generic_type of pdr_cfg : constant is 1;
    attribute mti_svvh_generic_type of ndr_cfg : constant is 1;
    attribute mti_svvh_generic_type of keep_cfg : constant is 1;
    attribute mti_svvh_generic_type of term_pu_en : constant is 1;
    attribute mti_svvh_generic_type of term_pd_en : constant is 1;
    attribute mti_svvh_generic_type of rx_dig_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of rx_hstl_sstl_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of tpd_cfg : constant is 1;
    attribute mti_svvh_generic_type of tpu_cfg : constant is 1;
    attribute mti_svvh_generic_type of cfg_trm : constant is 1;
    attribute mti_svvh_generic_type of cfg_trm_sel : constant is 1;
    attribute mti_svvh_generic_type of in_del : constant is 1;
    attribute mti_svvh_generic_type of out_del : constant is 1;
    attribute mti_svvh_generic_type of cfg_test_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_userio_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_use_cal0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_gsclk_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_gsclk90_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_gsclk180_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_gsclk270_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_gate_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_gate_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_rstn_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_rstn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_setn_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_setn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_setn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_setn_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_ddr : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_dqs : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd0_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd1_inv : constant is 1;
    attribute mti_svvh_generic_type of cfg_d_en : constant is 1;
    attribute mti_svvh_generic_type of cfg_clkout_sel : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_out : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_sel : constant is 1;
end M7A_IO_DDRSG;
