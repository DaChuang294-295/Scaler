library verilog;
use verilog.vl_types.all;
entity VCC is
    port(
        Y               : out    vl_logic
    );
end VCC;
