.box 1 demo_sd_to_lcd_ipc_adder_8 17 9
.input 1 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7]
.output 1 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] CO
.delay 1
-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	
400	300	200	-	-	-	-	-	400	400	300	200	100	-	-	-	-	
500	400	300	200	-	-	-	-	500	500	400	300	200	100	-	-	-	
600	500	400	300	200	-	-	-	600	600	500	400	300	200	100	-	-	
700	600	500	400	300	200	-	-	700	700	600	500	400	300	200	100	-	
800	700	600	500	400	300	200	-	800	800	700	600	500	400	300	200	100	
900	800	700	600	500	400	300	200	900	900	800	700	600	500	400	300	200	


