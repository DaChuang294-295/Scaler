library verilog;
use verilog.vl_types.all;
entity M7S_IO_LVDS is
    generic(
        cfg_nc          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ldr_cfg         : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_lvds_en_cfg  : vl_logic := Hi0;
        term_diff_en_cfg: vl_logic := Hi0;
        lvds_tx_en_cfg  : vl_logic := Hi0;
        cml_tx_en_cfg   : vl_logic := Hi0;
        td_cfg          : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        cfg_gear_mode48 : vl_logic := Hi0;
        cfg_gear_mode7  : vl_logic := Hi0;
        cfg_algn_rsn_sel: vl_logic := Hi0;
        ns_lv_fastestn_1: vl_logic := Hi0;
        cfg_userio_en_1 : vl_logic := Hi0;
        cfg_sclk_inv_1  : vl_logic := Hi0;
        cfg_sclk_gate_sel_1: vl_logic := Hi0;
        cfg_eclk_gate_sel_1: vl_logic := Hi0;
        cfg_eclk90_gate_sel_1: vl_logic := Hi0;
        cfg_sclk_en_1   : vl_logic := Hi0;
        cfg_fclk_en_1   : vl_logic := Hi0;
        cfg_eclk_en_1   : vl_logic := Hi0;
        cfg_eclk90_en_1 : vl_logic := Hi0;
        cfg_rstn_inv_1  : vl_logic := Hi0;
        cfg_oen_rstn_en_1: vl_logic := Hi0;
        cfg_od_rstn_en_1: vl_logic := Hi0;
        cfg_id_rstn_en_1: vl_logic := Hi0;
        cfg_setn_inv_1  : vl_logic := Hi0;
        cfg_oen_setn_en_1: vl_logic := Hi0;
        cfg_od_setn_en_1: vl_logic := Hi0;
        cfg_id_setn_en_1: vl_logic := Hi0;
        cfg_txd0_inv_1  : vl_logic := Hi0;
        cfg_txd1_inv_1  : vl_logic := Hi0;
        cfg_txd2_inv_1  : vl_logic := Hi0;
        cfg_txd3_inv_1  : vl_logic := Hi0;
        cfg_d_en_1      : vl_logic := Hi0;
        cfg_sclk_out_1  : vl_logic := Hi0;
        cfg_clkout_sel_1: vl_logic := Hi0;
        cfg_od_sel_1    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_oen_inv_1   : vl_logic := Hi0;
        cfg_oen_sel_1   : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_gear_1      : vl_logic := Hi0;
        cfg_slave_en_1  : vl_logic := Hi0;
        cfg_id_sel_1    : vl_logic := Hi0;
        ns_lv_cfg_1     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pdr_cfg_1       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ndr_cfg_1       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_dig_en_cfg_1 : vl_logic := Hi0;
        keep_cfg_1      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        in_del_1        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        out_del_1       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ns_lv_fastestn_0: vl_logic := Hi0;
        cfg_userio_en_0 : vl_logic := Hi0;
        cfg_sclk_inv_0  : vl_logic := Hi0;
        cfg_sclk_gate_sel_0: vl_logic := Hi0;
        cfg_eclk_gate_sel_0: vl_logic := Hi0;
        cfg_eclk90_gate_sel_0: vl_logic := Hi0;
        cfg_sclk_en_0   : vl_logic := Hi0;
        cfg_fclk_en_0   : vl_logic := Hi0;
        cfg_eclk_en_0   : vl_logic := Hi0;
        cfg_eclk90_en_0 : vl_logic := Hi0;
        cfg_rstn_inv_0  : vl_logic := Hi0;
        cfg_oen_rstn_en_0: vl_logic := Hi0;
        cfg_od_rstn_en_0: vl_logic := Hi0;
        cfg_id_rstn_en_0: vl_logic := Hi0;
        cfg_setn_inv_0  : vl_logic := Hi0;
        cfg_oen_setn_en_0: vl_logic := Hi0;
        cfg_od_setn_en_0: vl_logic := Hi0;
        cfg_id_setn_en_0: vl_logic := Hi0;
        cfg_txd0_inv_0  : vl_logic := Hi0;
        cfg_txd1_inv_0  : vl_logic := Hi0;
        cfg_txd2_inv_0  : vl_logic := Hi0;
        cfg_txd3_inv_0  : vl_logic := Hi0;
        cfg_d_en_0      : vl_logic := Hi0;
        cfg_sclk_out_0  : vl_logic := Hi0;
        cfg_clkout_sel_0: vl_logic := Hi0;
        cfg_od_sel_0    : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_oen_inv_0   : vl_logic := Hi0;
        cfg_oen_sel_0   : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        cfg_gear_0      : vl_logic := Hi0;
        cfg_slave_en_0  : vl_logic := Hi0;
        cfg_id_sel_0    : vl_logic := Hi0;
        ns_lv_cfg_0     : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        pdr_cfg_0       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        ndr_cfg_0       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        rx_dig_en_cfg_0 : vl_logic := Hi0;
        keep_cfg_0      : vl_logic_vector(0 to 1) := (Hi0, Hi0);
        in_del_0        : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        out_del_0       : vl_logic_vector(0 to 3) := (Hi0, Hi0, Hi0, Hi0);
        optional_function: string  := ""
    );
    port(
        id_1            : out    vl_logic;
        id_0            : out    vl_logic;
        id_q_1          : out    vl_logic_vector(3 downto 0);
        id_q_0          : out    vl_logic_vector(3 downto 0);
        align_rstn      : in     vl_logic;
        alignwd         : in     vl_logic;
        clk_en_1        : in     vl_logic;
        clk_en_0        : in     vl_logic;
        io_reg_clk      : out    vl_logic;
        geclk           : in     vl_logic;
        geclk90         : in     vl_logic;
        geclk180        : in     vl_logic;
        geclk270        : in     vl_logic;
        od_d_1          : in     vl_logic_vector(3 downto 0);
        od_d_0          : in     vl_logic_vector(3 downto 0);
        oen_1           : in     vl_logic;
        oen_0           : in     vl_logic;
        clk_0           : in     vl_logic;
        clk_1           : in     vl_logic;
        rstn_0          : in     vl_logic;
        rstn_1          : in     vl_logic;
        setn_0          : in     vl_logic;
        setn_1          : in     vl_logic;
        PAD1            : inout  vl_logic;
        PAD0            : inout  vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of cfg_nc : constant is 1;
    attribute mti_svvh_generic_type of ldr_cfg : constant is 1;
    attribute mti_svvh_generic_type of rx_lvds_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of term_diff_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of lvds_tx_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of cml_tx_en_cfg : constant is 1;
    attribute mti_svvh_generic_type of td_cfg : constant is 1;
    attribute mti_svvh_generic_type of cfg_gear_mode48 : constant is 1;
    attribute mti_svvh_generic_type of cfg_gear_mode7 : constant is 1;
    attribute mti_svvh_generic_type of cfg_algn_rsn_sel : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_fastestn_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_userio_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_gate_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk_gate_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk90_gate_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk90_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_rstn_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_rstn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_rstn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_rstn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_setn_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_setn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_setn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_setn_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd0_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd1_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd2_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd3_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_d_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_out_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_clkout_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_inv_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_gear_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_slave_en_1 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_sel_1 : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_cfg_1 : constant is 1;
    attribute mti_svvh_generic_type of pdr_cfg_1 : constant is 1;
    attribute mti_svvh_generic_type of ndr_cfg_1 : constant is 1;
    attribute mti_svvh_generic_type of rx_dig_en_cfg_1 : constant is 1;
    attribute mti_svvh_generic_type of keep_cfg_1 : constant is 1;
    attribute mti_svvh_generic_type of in_del_1 : constant is 1;
    attribute mti_svvh_generic_type of out_del_1 : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_fastestn_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_userio_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_gate_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk_gate_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk90_gate_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_fclk_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_eclk90_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_rstn_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_rstn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_rstn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_rstn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_setn_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_setn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_setn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_setn_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd0_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd1_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd2_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_txd3_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_d_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_sclk_out_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_clkout_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_od_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_inv_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_oen_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_gear_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_slave_en_0 : constant is 1;
    attribute mti_svvh_generic_type of cfg_id_sel_0 : constant is 1;
    attribute mti_svvh_generic_type of ns_lv_cfg_0 : constant is 1;
    attribute mti_svvh_generic_type of pdr_cfg_0 : constant is 1;
    attribute mti_svvh_generic_type of ndr_cfg_0 : constant is 1;
    attribute mti_svvh_generic_type of rx_dig_en_cfg_0 : constant is 1;
    attribute mti_svvh_generic_type of keep_cfg_0 : constant is 1;
    attribute mti_svvh_generic_type of in_del_0 : constant is 1;
    attribute mti_svvh_generic_type of out_del_0 : constant is 1;
    attribute mti_svvh_generic_type of optional_function : constant is 1;
end M7S_IO_LVDS;
