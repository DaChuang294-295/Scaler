module scaler_ipc_adder_11(CA, CI, CO, DX, SUM);
  input [10:0] CA;
  input CI;
  output CO;
  input [10:0] DX;
  output [10:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(CO), 
        .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_12(CA, CI, CO, DX, SUM);
  input [11:0] CA;
  input CI;
  output CO;
  input [11:0] DX;
  output [11:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(CO), 
        .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_14(CA, CI, CO, DX, SUM);
  input [13:0] CA;
  input CI;
  output CO;
  input [13:0] DX;
  output [13:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(CO), 
        .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_17(CA, CI, CO, DX, SUM);
  input [16:0] CA;
  input CI;
  output CO;
  input [16:0] DX;
  output [16:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(CO), 
        .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_18(CA, CI, CO, DX, SUM);
  input [17:0] CA;
  input CI;
  output CO;
  input [17:0] DX;
  output [17:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_16|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(
        \MUXCO_16|COUT_net ), .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_17 ( .AIN(CA[17]), .CIN(\MUXCO_16|COUT_net ), .COUT(CO), 
        .CSEL(DX[17]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_17 ( .CIN(\MUXCO_16|COUT_net ), .DIN(DX[17]), .SUM(
        SUM[17]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_34(CA, CI, CO, DX, SUM);
  input [33:0] CA;
  input CI;
  output CO;
  input [33:0] DX;
  output [33:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_16|COUT_net ;
    wire \MUXCO_17|COUT_net ;
    wire \MUXCO_18|COUT_net ;
    wire \MUXCO_19|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_20|COUT_net ;
    wire \MUXCO_21|COUT_net ;
    wire \MUXCO_22|COUT_net ;
    wire \MUXCO_23|COUT_net ;
    wire \MUXCO_24|COUT_net ;
    wire \MUXCO_25|COUT_net ;
    wire \MUXCO_26|COUT_net ;
    wire \MUXCO_27|COUT_net ;
    wire \MUXCO_28|COUT_net ;
    wire \MUXCO_29|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_30|COUT_net ;
    wire \MUXCO_31|COUT_net ;
    wire \MUXCO_32|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(
        \MUXCO_16|COUT_net ), .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_17 ( .AIN(CA[17]), .CIN(\MUXCO_16|COUT_net ), .COUT(
        \MUXCO_17|COUT_net ), .CSEL(DX[17]) );
    CS_MUXCO_PRIM MUXCO_18 ( .AIN(CA[18]), .CIN(\MUXCO_17|COUT_net ), .COUT(
        \MUXCO_18|COUT_net ), .CSEL(DX[18]) );
    CS_MUXCO_PRIM MUXCO_19 ( .AIN(CA[19]), .CIN(\MUXCO_18|COUT_net ), .COUT(
        \MUXCO_19|COUT_net ), .CSEL(DX[19]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_20 ( .AIN(CA[20]), .CIN(\MUXCO_19|COUT_net ), .COUT(
        \MUXCO_20|COUT_net ), .CSEL(DX[20]) );
    CS_MUXCO_PRIM MUXCO_21 ( .AIN(CA[21]), .CIN(\MUXCO_20|COUT_net ), .COUT(
        \MUXCO_21|COUT_net ), .CSEL(DX[21]) );
    CS_MUXCO_PRIM MUXCO_22 ( .AIN(CA[22]), .CIN(\MUXCO_21|COUT_net ), .COUT(
        \MUXCO_22|COUT_net ), .CSEL(DX[22]) );
    CS_MUXCO_PRIM MUXCO_23 ( .AIN(CA[23]), .CIN(\MUXCO_22|COUT_net ), .COUT(
        \MUXCO_23|COUT_net ), .CSEL(DX[23]) );
    CS_MUXCO_PRIM MUXCO_24 ( .AIN(CA[24]), .CIN(\MUXCO_23|COUT_net ), .COUT(
        \MUXCO_24|COUT_net ), .CSEL(DX[24]) );
    CS_MUXCO_PRIM MUXCO_25 ( .AIN(CA[25]), .CIN(\MUXCO_24|COUT_net ), .COUT(
        \MUXCO_25|COUT_net ), .CSEL(DX[25]) );
    CS_MUXCO_PRIM MUXCO_26 ( .AIN(CA[26]), .CIN(\MUXCO_25|COUT_net ), .COUT(
        \MUXCO_26|COUT_net ), .CSEL(DX[26]) );
    CS_MUXCO_PRIM MUXCO_27 ( .AIN(CA[27]), .CIN(\MUXCO_26|COUT_net ), .COUT(
        \MUXCO_27|COUT_net ), .CSEL(DX[27]) );
    CS_MUXCO_PRIM MUXCO_28 ( .AIN(CA[28]), .CIN(\MUXCO_27|COUT_net ), .COUT(
        \MUXCO_28|COUT_net ), .CSEL(DX[28]) );
    CS_MUXCO_PRIM MUXCO_29 ( .AIN(CA[29]), .CIN(\MUXCO_28|COUT_net ), .COUT(
        \MUXCO_29|COUT_net ), .CSEL(DX[29]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_30 ( .AIN(CA[30]), .CIN(\MUXCO_29|COUT_net ), .COUT(
        \MUXCO_30|COUT_net ), .CSEL(DX[30]) );
    CS_MUXCO_PRIM MUXCO_31 ( .AIN(CA[31]), .CIN(\MUXCO_30|COUT_net ), .COUT(
        \MUXCO_31|COUT_net ), .CSEL(DX[31]) );
    CS_MUXCO_PRIM MUXCO_32 ( .AIN(CA[32]), .CIN(\MUXCO_31|COUT_net ), .COUT(
        \MUXCO_32|COUT_net ), .CSEL(DX[32]) );
    CS_MUXCO_PRIM MUXCO_33 ( .AIN(CA[33]), .CIN(\MUXCO_32|COUT_net ), .COUT(CO), 
        .CSEL(DX[33]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_17 ( .CIN(\MUXCO_16|COUT_net ), .DIN(DX[17]), .SUM(
        SUM[17]) );
    CS_XORCI_PRIM XORCI_18 ( .CIN(\MUXCO_17|COUT_net ), .DIN(DX[18]), .SUM(
        SUM[18]) );
    CS_XORCI_PRIM XORCI_19 ( .CIN(\MUXCO_18|COUT_net ), .DIN(DX[19]), .SUM(
        SUM[19]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_20 ( .CIN(\MUXCO_19|COUT_net ), .DIN(DX[20]), .SUM(
        SUM[20]) );
    CS_XORCI_PRIM XORCI_21 ( .CIN(\MUXCO_20|COUT_net ), .DIN(DX[21]), .SUM(
        SUM[21]) );
    CS_XORCI_PRIM XORCI_22 ( .CIN(\MUXCO_21|COUT_net ), .DIN(DX[22]), .SUM(
        SUM[22]) );
    CS_XORCI_PRIM XORCI_23 ( .CIN(\MUXCO_22|COUT_net ), .DIN(DX[23]), .SUM(
        SUM[23]) );
    CS_XORCI_PRIM XORCI_24 ( .CIN(\MUXCO_23|COUT_net ), .DIN(DX[24]), .SUM(
        SUM[24]) );
    CS_XORCI_PRIM XORCI_25 ( .CIN(\MUXCO_24|COUT_net ), .DIN(DX[25]), .SUM(
        SUM[25]) );
    CS_XORCI_PRIM XORCI_26 ( .CIN(\MUXCO_25|COUT_net ), .DIN(DX[26]), .SUM(
        SUM[26]) );
    CS_XORCI_PRIM XORCI_27 ( .CIN(\MUXCO_26|COUT_net ), .DIN(DX[27]), .SUM(
        SUM[27]) );
    CS_XORCI_PRIM XORCI_28 ( .CIN(\MUXCO_27|COUT_net ), .DIN(DX[28]), .SUM(
        SUM[28]) );
    CS_XORCI_PRIM XORCI_29 ( .CIN(\MUXCO_28|COUT_net ), .DIN(DX[29]), .SUM(
        SUM[29]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_30 ( .CIN(\MUXCO_29|COUT_net ), .DIN(DX[30]), .SUM(
        SUM[30]) );
    CS_XORCI_PRIM XORCI_31 ( .CIN(\MUXCO_30|COUT_net ), .DIN(DX[31]), .SUM(
        SUM[31]) );
    CS_XORCI_PRIM XORCI_32 ( .CIN(\MUXCO_31|COUT_net ), .DIN(DX[32]), .SUM(
        SUM[32]) );
    CS_XORCI_PRIM XORCI_33 ( .CIN(\MUXCO_32|COUT_net ), .DIN(DX[33]), .SUM(
        SUM[33]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_7(CA, CI, CO, DX, SUM);
  input [6:0] CA;
  input CI;
  output CO;
  input [6:0] DX;
  output [6:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(CO), 
        .CSEL(DX[6]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
endmodule


module scaler_ipc_adder_8(CA, CI, CO, DX, SUM);
  input [7:0] CA;
  input CI;
  output CO;
  input [7:0] DX;
  output [7:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(CO), 
        .CSEL(DX[7]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
endmodule


module scaler ( HS, VS, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u135_mac, a_acc_en_cal1_u136_mac,
           a_acc_en_cal1_u137_mac, a_acc_en_cal1_u138_mac, a_acc_en_cal1_u139_mac,
           a_acc_en_cal1_u140_mac, a_acc_en_cal1_u141_mac, a_acc_en_cal1_u142_mac,
           a_acc_en_cal1_u143_mac, a_acc_en_cal1_u144_mac, a_acc_en_cal1_u145_mac,
           a_acc_en_cal1_u146_mac, a_acc_en_coefcal1_u63_mac, a_acc_en_coefcal1_u64_mac,
           a_acc_en_coefcal1_u64_mac_0_, \a_dinx[0]_cal1_u134_mac , \a_dinx[0]_cal1_u135_mac ,
           \a_dinx[0]_cal1_u136_mac , \a_dinx[0]_cal1_u137_mac , \a_dinx[0]_cal1_u138_mac ,
           \a_dinx[0]_cal1_u139_mac , \a_dinx[0]_cal1_u140_mac , \a_dinx[0]_cal1_u141_mac ,
           \a_dinx[0]_cal1_u142_mac , \a_dinx[0]_cal1_u143_mac , \a_dinx[0]_cal1_u144_mac ,
           \a_dinx[0]_cal1_u145_mac , \a_dinx[0]_cal1_u146_mac , \a_dinx[0]_coefcal1_u63_mac ,
           \a_dinx[0]_coefcal1_u64_mac , \a_dinx[0]_coefcal1_u64_mac_0_ ,
           \a_dinx[10]_cal1_u134_mac , \a_dinx[10]_cal1_u135_mac , \a_dinx[10]_cal1_u136_mac ,
           \a_dinx[10]_cal1_u137_mac , \a_dinx[10]_cal1_u138_mac , \a_dinx[10]_cal1_u139_mac ,
           \a_dinx[10]_cal1_u140_mac , \a_dinx[10]_cal1_u141_mac , \a_dinx[10]_cal1_u142_mac ,
           \a_dinx[10]_cal1_u143_mac , \a_dinx[10]_cal1_u144_mac , \a_dinx[10]_cal1_u145_mac ,
           \a_dinx[10]_cal1_u146_mac , \a_dinx[10]_coefcal1_u63_mac , \a_dinx[10]_coefcal1_u64_mac ,
           \a_dinx[10]_coefcal1_u64_mac_0_ , \a_dinx[11]_cal1_u134_mac , \a_dinx[11]_cal1_u135_mac ,
           \a_dinx[11]_cal1_u136_mac , \a_dinx[11]_cal1_u137_mac , \a_dinx[11]_cal1_u138_mac ,
           \a_dinx[11]_cal1_u139_mac , \a_dinx[11]_cal1_u140_mac , \a_dinx[11]_cal1_u141_mac ,
           \a_dinx[11]_cal1_u142_mac , \a_dinx[11]_cal1_u143_mac , \a_dinx[11]_cal1_u144_mac ,
           \a_dinx[11]_cal1_u145_mac , \a_dinx[11]_cal1_u146_mac , \a_dinx[11]_coefcal1_u63_mac ,
           \a_dinx[11]_coefcal1_u64_mac , \a_dinx[11]_coefcal1_u64_mac_0_ ,
           \a_dinx[12]_cal1_u134_mac , \a_dinx[12]_cal1_u135_mac , \a_dinx[12]_cal1_u136_mac ,
           \a_dinx[12]_cal1_u137_mac , \a_dinx[12]_cal1_u138_mac , \a_dinx[12]_cal1_u139_mac ,
           \a_dinx[12]_cal1_u140_mac , \a_dinx[12]_cal1_u141_mac , \a_dinx[12]_cal1_u142_mac ,
           \a_dinx[12]_cal1_u143_mac , \a_dinx[12]_cal1_u144_mac , \a_dinx[12]_cal1_u145_mac ,
           \a_dinx[12]_cal1_u146_mac , \a_dinx[12]_coefcal1_u63_mac , \a_dinx[12]_coefcal1_u64_mac ,
           \a_dinx[12]_coefcal1_u64_mac_0_ , \a_dinx[13]_cal1_u134_mac , \a_dinx[13]_cal1_u135_mac ,
           \a_dinx[13]_cal1_u136_mac , \a_dinx[13]_cal1_u137_mac , \a_dinx[13]_cal1_u138_mac ,
           \a_dinx[13]_cal1_u139_mac , \a_dinx[13]_cal1_u140_mac , \a_dinx[13]_cal1_u141_mac ,
           \a_dinx[13]_cal1_u142_mac , \a_dinx[13]_cal1_u143_mac , \a_dinx[13]_cal1_u144_mac ,
           \a_dinx[13]_cal1_u145_mac , \a_dinx[13]_cal1_u146_mac , \a_dinx[13]_coefcal1_u63_mac ,
           \a_dinx[13]_coefcal1_u64_mac , \a_dinx[13]_coefcal1_u64_mac_0_ ,
           \a_dinx[1]_cal1_u134_mac , \a_dinx[1]_cal1_u135_mac , \a_dinx[1]_cal1_u136_mac ,
           \a_dinx[1]_cal1_u137_mac , \a_dinx[1]_cal1_u138_mac , \a_dinx[1]_cal1_u139_mac ,
           \a_dinx[1]_cal1_u140_mac , \a_dinx[1]_cal1_u141_mac , \a_dinx[1]_cal1_u142_mac ,
           \a_dinx[1]_cal1_u143_mac , \a_dinx[1]_cal1_u144_mac , \a_dinx[1]_cal1_u145_mac ,
           \a_dinx[1]_cal1_u146_mac , \a_dinx[1]_coefcal1_u63_mac , \a_dinx[1]_coefcal1_u64_mac ,
           \a_dinx[1]_coefcal1_u64_mac_0_ , \a_dinx[2]_cal1_u134_mac , \a_dinx[2]_cal1_u135_mac ,
           \a_dinx[2]_cal1_u136_mac , \a_dinx[2]_cal1_u137_mac , \a_dinx[2]_cal1_u138_mac ,
           \a_dinx[2]_cal1_u139_mac , \a_dinx[2]_cal1_u140_mac , \a_dinx[2]_cal1_u141_mac ,
           \a_dinx[2]_cal1_u142_mac , \a_dinx[2]_cal1_u143_mac , \a_dinx[2]_cal1_u144_mac ,
           \a_dinx[2]_cal1_u145_mac , \a_dinx[2]_cal1_u146_mac , \a_dinx[2]_coefcal1_u63_mac ,
           \a_dinx[2]_coefcal1_u64_mac , \a_dinx[2]_coefcal1_u64_mac_0_ ,
           \a_dinx[3]_cal1_u134_mac , \a_dinx[3]_cal1_u135_mac , \a_dinx[3]_cal1_u136_mac ,
           \a_dinx[3]_cal1_u137_mac , \a_dinx[3]_cal1_u138_mac , \a_dinx[3]_cal1_u139_mac ,
           \a_dinx[3]_cal1_u140_mac , \a_dinx[3]_cal1_u141_mac , \a_dinx[3]_cal1_u142_mac ,
           \a_dinx[3]_cal1_u143_mac , \a_dinx[3]_cal1_u144_mac , \a_dinx[3]_cal1_u145_mac ,
           \a_dinx[3]_cal1_u146_mac , \a_dinx[3]_coefcal1_u63_mac , \a_dinx[3]_coefcal1_u64_mac ,
           \a_dinx[3]_coefcal1_u64_mac_0_ , \a_dinx[4]_cal1_u134_mac , \a_dinx[4]_cal1_u135_mac ,
           \a_dinx[4]_cal1_u136_mac , \a_dinx[4]_cal1_u137_mac , \a_dinx[4]_cal1_u138_mac ,
           \a_dinx[4]_cal1_u139_mac , \a_dinx[4]_cal1_u140_mac , \a_dinx[4]_cal1_u141_mac ,
           \a_dinx[4]_cal1_u142_mac , \a_dinx[4]_cal1_u143_mac , \a_dinx[4]_cal1_u144_mac ,
           \a_dinx[4]_cal1_u145_mac , \a_dinx[4]_cal1_u146_mac , \a_dinx[4]_coefcal1_u63_mac ,
           \a_dinx[4]_coefcal1_u64_mac , \a_dinx[4]_coefcal1_u64_mac_0_ ,
           \a_dinx[5]_cal1_u134_mac , \a_dinx[5]_cal1_u135_mac , \a_dinx[5]_cal1_u136_mac ,
           \a_dinx[5]_cal1_u137_mac , \a_dinx[5]_cal1_u138_mac , \a_dinx[5]_cal1_u139_mac ,
           \a_dinx[5]_cal1_u140_mac , \a_dinx[5]_cal1_u141_mac , \a_dinx[5]_cal1_u142_mac ,
           \a_dinx[5]_cal1_u143_mac , \a_dinx[5]_cal1_u144_mac , \a_dinx[5]_cal1_u145_mac ,
           \a_dinx[5]_cal1_u146_mac , \a_dinx[5]_coefcal1_u63_mac , \a_dinx[5]_coefcal1_u64_mac ,
           \a_dinx[5]_coefcal1_u64_mac_0_ , \a_dinx[6]_cal1_u134_mac , \a_dinx[6]_cal1_u135_mac ,
           \a_dinx[6]_cal1_u136_mac , \a_dinx[6]_cal1_u137_mac , \a_dinx[6]_cal1_u138_mac ,
           \a_dinx[6]_cal1_u139_mac , \a_dinx[6]_cal1_u140_mac , \a_dinx[6]_cal1_u141_mac ,
           \a_dinx[6]_cal1_u142_mac , \a_dinx[6]_cal1_u143_mac , \a_dinx[6]_cal1_u144_mac ,
           \a_dinx[6]_cal1_u145_mac , \a_dinx[6]_cal1_u146_mac , \a_dinx[6]_coefcal1_u63_mac ,
           \a_dinx[6]_coefcal1_u64_mac , \a_dinx[6]_coefcal1_u64_mac_0_ ,
           \a_dinx[7]_cal1_u134_mac , \a_dinx[7]_cal1_u135_mac , \a_dinx[7]_cal1_u136_mac ,
           \a_dinx[7]_cal1_u137_mac , \a_dinx[7]_cal1_u138_mac , \a_dinx[7]_cal1_u139_mac ,
           \a_dinx[7]_cal1_u140_mac , \a_dinx[7]_cal1_u141_mac , \a_dinx[7]_cal1_u142_mac ,
           \a_dinx[7]_cal1_u143_mac , \a_dinx[7]_cal1_u144_mac , \a_dinx[7]_cal1_u145_mac ,
           \a_dinx[7]_cal1_u146_mac , \a_dinx[7]_coefcal1_u63_mac , \a_dinx[7]_coefcal1_u64_mac ,
           \a_dinx[7]_coefcal1_u64_mac_0_ , \a_dinx[8]_cal1_u134_mac , \a_dinx[8]_cal1_u135_mac ,
           \a_dinx[8]_cal1_u136_mac , \a_dinx[8]_cal1_u137_mac , \a_dinx[8]_cal1_u138_mac ,
           \a_dinx[8]_cal1_u139_mac , \a_dinx[8]_cal1_u140_mac , \a_dinx[8]_cal1_u141_mac ,
           \a_dinx[8]_cal1_u142_mac , \a_dinx[8]_cal1_u143_mac , \a_dinx[8]_cal1_u144_mac ,
           \a_dinx[8]_cal1_u145_mac , \a_dinx[8]_cal1_u146_mac , \a_dinx[8]_coefcal1_u63_mac ,
           \a_dinx[8]_coefcal1_u64_mac , \a_dinx[8]_coefcal1_u64_mac_0_ ,
           \a_dinx[9]_cal1_u134_mac , \a_dinx[9]_cal1_u135_mac , \a_dinx[9]_cal1_u136_mac ,
           \a_dinx[9]_cal1_u137_mac , \a_dinx[9]_cal1_u138_mac , \a_dinx[9]_cal1_u139_mac ,
           \a_dinx[9]_cal1_u140_mac , \a_dinx[9]_cal1_u141_mac , \a_dinx[9]_cal1_u142_mac ,
           \a_dinx[9]_cal1_u143_mac , \a_dinx[9]_cal1_u144_mac , \a_dinx[9]_cal1_u145_mac ,
           \a_dinx[9]_cal1_u146_mac , \a_dinx[9]_coefcal1_u63_mac , \a_dinx[9]_coefcal1_u64_mac ,
           \a_dinx[9]_coefcal1_u64_mac_0_ , a_dinxy_cen_cal1_u134_mac, a_dinxy_cen_cal1_u135_mac,
           a_dinxy_cen_cal1_u136_mac, a_dinxy_cen_cal1_u137_mac, a_dinxy_cen_cal1_u138_mac,
           a_dinxy_cen_cal1_u139_mac, a_dinxy_cen_cal1_u140_mac, a_dinxy_cen_cal1_u141_mac,
           a_dinxy_cen_cal1_u142_mac, a_dinxy_cen_cal1_u143_mac, a_dinxy_cen_cal1_u144_mac,
           a_dinxy_cen_cal1_u145_mac, a_dinxy_cen_cal1_u146_mac, a_dinxy_cen_coefcal1_u63_mac,
           a_dinxy_cen_coefcal1_u64_mac, a_dinxy_cen_coefcal1_u64_mac_0_,
           \a_diny[0]_cal1_u134_mac , \a_diny[0]_cal1_u135_mac , \a_diny[0]_cal1_u136_mac ,
           \a_diny[0]_cal1_u137_mac , \a_diny[0]_cal1_u138_mac , \a_diny[0]_cal1_u139_mac ,
           \a_diny[0]_cal1_u140_mac , \a_diny[0]_cal1_u141_mac , \a_diny[0]_cal1_u142_mac ,
           \a_diny[0]_cal1_u143_mac , \a_diny[0]_cal1_u144_mac , \a_diny[0]_cal1_u145_mac ,
           \a_diny[0]_cal1_u146_mac , \a_diny[0]_coefcal1_u63_mac , \a_diny[0]_coefcal1_u64_mac ,
           \a_diny[0]_coefcal1_u64_mac_0_ , \a_diny[1]_cal1_u134_mac , \a_diny[1]_cal1_u135_mac ,
           \a_diny[1]_cal1_u136_mac , \a_diny[1]_cal1_u137_mac , \a_diny[1]_cal1_u138_mac ,
           \a_diny[1]_cal1_u139_mac , \a_diny[1]_cal1_u140_mac , \a_diny[1]_cal1_u141_mac ,
           \a_diny[1]_cal1_u142_mac , \a_diny[1]_cal1_u143_mac , \a_diny[1]_cal1_u144_mac ,
           \a_diny[1]_cal1_u145_mac , \a_diny[1]_cal1_u146_mac , \a_diny[1]_coefcal1_u63_mac ,
           \a_diny[1]_coefcal1_u64_mac , \a_diny[1]_coefcal1_u64_mac_0_ ,
           \a_diny[2]_cal1_u134_mac , \a_diny[2]_cal1_u135_mac , \a_diny[2]_cal1_u136_mac ,
           \a_diny[2]_cal1_u137_mac , \a_diny[2]_cal1_u138_mac , \a_diny[2]_cal1_u139_mac ,
           \a_diny[2]_cal1_u140_mac , \a_diny[2]_cal1_u141_mac , \a_diny[2]_cal1_u142_mac ,
           \a_diny[2]_cal1_u143_mac , \a_diny[2]_cal1_u144_mac , \a_diny[2]_cal1_u145_mac ,
           \a_diny[2]_cal1_u146_mac , \a_diny[2]_coefcal1_u63_mac , \a_diny[2]_coefcal1_u64_mac ,
           \a_diny[2]_coefcal1_u64_mac_0_ , \a_diny[3]_cal1_u134_mac , \a_diny[3]_cal1_u135_mac ,
           \a_diny[3]_cal1_u136_mac , \a_diny[3]_cal1_u137_mac , \a_diny[3]_cal1_u138_mac ,
           \a_diny[3]_cal1_u139_mac , \a_diny[3]_cal1_u140_mac , \a_diny[3]_cal1_u141_mac ,
           \a_diny[3]_cal1_u142_mac , \a_diny[3]_cal1_u143_mac , \a_diny[3]_cal1_u144_mac ,
           \a_diny[3]_cal1_u145_mac , \a_diny[3]_cal1_u146_mac , \a_diny[3]_coefcal1_u63_mac ,
           \a_diny[3]_coefcal1_u64_mac , \a_diny[3]_coefcal1_u64_mac_0_ ,
           \a_diny[4]_cal1_u134_mac , \a_diny[4]_cal1_u135_mac , \a_diny[4]_cal1_u136_mac ,
           \a_diny[4]_cal1_u137_mac , \a_diny[4]_cal1_u138_mac , \a_diny[4]_cal1_u139_mac ,
           \a_diny[4]_cal1_u140_mac , \a_diny[4]_cal1_u141_mac , \a_diny[4]_cal1_u142_mac ,
           \a_diny[4]_cal1_u143_mac , \a_diny[4]_cal1_u144_mac , \a_diny[4]_cal1_u145_mac ,
           \a_diny[4]_cal1_u146_mac , \a_diny[4]_coefcal1_u63_mac , \a_diny[4]_coefcal1_u64_mac ,
           \a_diny[4]_coefcal1_u64_mac_0_ , \a_diny[5]_cal1_u134_mac , \a_diny[5]_cal1_u135_mac ,
           \a_diny[5]_cal1_u136_mac , \a_diny[5]_cal1_u137_mac , \a_diny[5]_cal1_u138_mac ,
           \a_diny[5]_cal1_u139_mac , \a_diny[5]_cal1_u140_mac , \a_diny[5]_cal1_u141_mac ,
           \a_diny[5]_cal1_u142_mac , \a_diny[5]_cal1_u143_mac , \a_diny[5]_cal1_u144_mac ,
           \a_diny[5]_cal1_u145_mac , \a_diny[5]_cal1_u146_mac , \a_diny[5]_coefcal1_u63_mac ,
           \a_diny[5]_coefcal1_u64_mac , \a_diny[5]_coefcal1_u64_mac_0_ ,
           \a_diny[6]_cal1_u134_mac , \a_diny[6]_cal1_u135_mac , \a_diny[6]_cal1_u136_mac ,
           \a_diny[6]_cal1_u137_mac , \a_diny[6]_cal1_u138_mac , \a_diny[6]_cal1_u139_mac ,
           \a_diny[6]_cal1_u140_mac , \a_diny[6]_cal1_u141_mac , \a_diny[6]_cal1_u142_mac ,
           \a_diny[6]_cal1_u143_mac , \a_diny[6]_cal1_u144_mac , \a_diny[6]_cal1_u145_mac ,
           \a_diny[6]_cal1_u146_mac , \a_diny[6]_coefcal1_u63_mac , \a_diny[6]_coefcal1_u64_mac ,
           \a_diny[6]_coefcal1_u64_mac_0_ , \a_diny[7]_cal1_u134_mac , \a_diny[7]_cal1_u135_mac ,
           \a_diny[7]_cal1_u136_mac , \a_diny[7]_cal1_u137_mac , \a_diny[7]_cal1_u138_mac ,
           \a_diny[7]_cal1_u139_mac , \a_diny[7]_cal1_u140_mac , \a_diny[7]_cal1_u141_mac ,
           \a_diny[7]_cal1_u142_mac , \a_diny[7]_cal1_u143_mac , \a_diny[7]_cal1_u144_mac ,
           \a_diny[7]_cal1_u145_mac , \a_diny[7]_cal1_u146_mac , \a_diny[7]_coefcal1_u63_mac ,
           \a_diny[7]_coefcal1_u64_mac , \a_diny[7]_coefcal1_u64_mac_0_ ,
           \a_diny[8]_cal1_u134_mac , \a_diny[8]_cal1_u135_mac , \a_diny[8]_cal1_u136_mac ,
           \a_diny[8]_cal1_u137_mac , \a_diny[8]_cal1_u138_mac , \a_diny[8]_cal1_u139_mac ,
           \a_diny[8]_cal1_u140_mac , \a_diny[8]_cal1_u141_mac , \a_diny[8]_cal1_u142_mac ,
           \a_diny[8]_cal1_u143_mac , \a_diny[8]_cal1_u144_mac , \a_diny[8]_cal1_u145_mac ,
           \a_diny[8]_cal1_u146_mac , \a_diny[8]_coefcal1_u63_mac , \a_diny[8]_coefcal1_u64_mac ,
           \a_diny[8]_coefcal1_u64_mac_0_ , \a_diny[9]_cal1_u134_mac , \a_diny[9]_cal1_u135_mac ,
           \a_diny[9]_cal1_u136_mac , \a_diny[9]_cal1_u137_mac , \a_diny[9]_cal1_u138_mac ,
           \a_diny[9]_cal1_u139_mac , \a_diny[9]_cal1_u140_mac , \a_diny[9]_cal1_u141_mac ,
           \a_diny[9]_cal1_u142_mac , \a_diny[9]_cal1_u143_mac , \a_diny[9]_cal1_u144_mac ,
           \a_diny[9]_cal1_u145_mac , \a_diny[9]_cal1_u146_mac , \a_diny[9]_coefcal1_u63_mac ,
           \a_diny[9]_coefcal1_u64_mac , \a_diny[9]_coefcal1_u64_mac_0_ ,
           a_dinz_cen_cal1_u134_mac, a_dinz_cen_cal1_u135_mac, a_dinz_cen_cal1_u136_mac,
           a_dinz_cen_cal1_u137_mac, a_dinz_cen_cal1_u138_mac, a_dinz_cen_cal1_u139_mac,
           a_dinz_cen_cal1_u140_mac, a_dinz_cen_cal1_u141_mac, a_dinz_cen_cal1_u142_mac,
           a_dinz_cen_cal1_u143_mac, a_dinz_cen_cal1_u144_mac, a_dinz_cen_cal1_u145_mac,
           a_dinz_cen_cal1_u146_mac, a_dinz_cen_coefcal1_u63_mac, a_dinz_cen_coefcal1_u64_mac,
           a_dinz_cen_coefcal1_u64_mac_0_, a_dinz_en_cal1_u134_mac, a_dinz_en_cal1_u135_mac,
           a_dinz_en_cal1_u136_mac, a_dinz_en_cal1_u137_mac, a_dinz_en_cal1_u138_mac,
           a_dinz_en_cal1_u139_mac, a_dinz_en_cal1_u140_mac, a_dinz_en_cal1_u141_mac,
           a_dinz_en_cal1_u142_mac, a_dinz_en_cal1_u143_mac, a_dinz_en_cal1_u144_mac,
           a_dinz_en_cal1_u145_mac, a_dinz_en_cal1_u146_mac, a_dinz_en_coefcal1_u63_mac,
           a_dinz_en_coefcal1_u64_mac, a_dinz_en_coefcal1_u64_mac_0_, a_in_sr_cal1_u134_mac,
           a_in_sr_cal1_u135_mac, a_in_sr_cal1_u136_mac, a_in_sr_cal1_u137_mac,
           a_in_sr_cal1_u138_mac, a_in_sr_cal1_u139_mac, a_in_sr_cal1_u140_mac,
           a_in_sr_cal1_u141_mac, a_in_sr_cal1_u142_mac, a_in_sr_cal1_u143_mac,
           a_in_sr_cal1_u144_mac, a_in_sr_cal1_u145_mac, a_in_sr_cal1_u146_mac,
           a_in_sr_coefcal1_u63_mac, a_in_sr_coefcal1_u64_mac, a_in_sr_coefcal1_u64_mac_0_,
           \a_mac_out[0]_coefcal1_u63_mac , \a_mac_out[0]_coefcal1_u64_mac ,
           \a_mac_out[0]_coefcal1_u64_mac_0_ , \a_mac_out[10]_cal1_u134_mac ,
           \a_mac_out[10]_cal1_u135_mac , \a_mac_out[10]_cal1_u136_mac , \a_mac_out[10]_cal1_u137_mac ,
           \a_mac_out[10]_cal1_u138_mac , \a_mac_out[10]_cal1_u139_mac , \a_mac_out[10]_cal1_u140_mac ,
           \a_mac_out[10]_cal1_u141_mac , \a_mac_out[10]_cal1_u142_mac , \a_mac_out[10]_cal1_u143_mac ,
           \a_mac_out[10]_cal1_u144_mac , \a_mac_out[10]_cal1_u145_mac , \a_mac_out[10]_cal1_u146_mac ,
           \a_mac_out[10]_coefcal1_u63_mac , \a_mac_out[10]_coefcal1_u64_mac ,
           \a_mac_out[10]_coefcal1_u64_mac_0_ , \a_mac_out[11]_cal1_u134_mac ,
           \a_mac_out[11]_cal1_u139_mac , \a_mac_out[11]_cal1_u140_mac , \a_mac_out[11]_cal1_u141_mac ,
           \a_mac_out[11]_cal1_u142_mac , \a_mac_out[11]_coefcal1_u63_mac ,
           \a_mac_out[11]_coefcal1_u64_mac , \a_mac_out[11]_coefcal1_u64_mac_0_ ,
           \a_mac_out[12]_coefcal1_u63_mac , \a_mac_out[12]_coefcal1_u64_mac ,
           \a_mac_out[12]_coefcal1_u64_mac_0_ , \a_mac_out[13]_coefcal1_u63_mac ,
           \a_mac_out[13]_coefcal1_u64_mac , \a_mac_out[14]_coefcal1_u63_mac ,
           \a_mac_out[14]_coefcal1_u64_mac , \a_mac_out[15]_coefcal1_u63_mac ,
           \a_mac_out[15]_coefcal1_u64_mac , \a_mac_out[16]_coefcal1_u63_mac ,
           \a_mac_out[16]_coefcal1_u64_mac , \a_mac_out[17]_coefcal1_u63_mac ,
           \a_mac_out[17]_coefcal1_u64_mac , \a_mac_out[18]_coefcal1_u63_mac ,
           \a_mac_out[18]_coefcal1_u64_mac , \a_mac_out[19]_coefcal1_u63_mac ,
           \a_mac_out[19]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u63_mac ,
           \a_mac_out[1]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u64_mac_0_ ,
           \a_mac_out[20]_coefcal1_u64_mac , \a_mac_out[21]_coefcal1_u64_mac ,
           \a_mac_out[22]_coefcal1_u64_mac , \a_mac_out[23]_coefcal1_u64_mac ,
           \a_mac_out[2]_coefcal1_u63_mac , \a_mac_out[2]_coefcal1_u64_mac ,
           \a_mac_out[2]_coefcal1_u64_mac_0_ , \a_mac_out[3]_coefcal1_u63_mac ,
           \a_mac_out[3]_coefcal1_u64_mac , \a_mac_out[3]_coefcal1_u64_mac_0_ ,
           \a_mac_out[4]_coefcal1_u63_mac , \a_mac_out[4]_coefcal1_u64_mac ,
           \a_mac_out[4]_coefcal1_u64_mac_0_ , \a_mac_out[5]_coefcal1_u63_mac ,
           \a_mac_out[5]_coefcal1_u64_mac , \a_mac_out[5]_coefcal1_u64_mac_0_ ,
           \a_mac_out[6]_cal1_u134_mac , \a_mac_out[6]_cal1_u135_mac , \a_mac_out[6]_cal1_u136_mac ,
           \a_mac_out[6]_cal1_u137_mac , \a_mac_out[6]_cal1_u138_mac , \a_mac_out[6]_cal1_u139_mac ,
           \a_mac_out[6]_cal1_u140_mac , \a_mac_out[6]_cal1_u141_mac , \a_mac_out[6]_cal1_u142_mac ,
           \a_mac_out[6]_cal1_u143_mac , \a_mac_out[6]_cal1_u144_mac , \a_mac_out[6]_cal1_u145_mac ,
           \a_mac_out[6]_cal1_u146_mac , \a_mac_out[6]_coefcal1_u63_mac ,
           \a_mac_out[6]_coefcal1_u64_mac , \a_mac_out[6]_coefcal1_u64_mac_0_ ,
           \a_mac_out[7]_cal1_u134_mac , \a_mac_out[7]_cal1_u135_mac , \a_mac_out[7]_cal1_u136_mac ,
           \a_mac_out[7]_cal1_u137_mac , \a_mac_out[7]_cal1_u138_mac , \a_mac_out[7]_cal1_u139_mac ,
           \a_mac_out[7]_cal1_u140_mac , \a_mac_out[7]_cal1_u141_mac , \a_mac_out[7]_cal1_u142_mac ,
           \a_mac_out[7]_cal1_u143_mac , \a_mac_out[7]_cal1_u144_mac , \a_mac_out[7]_cal1_u145_mac ,
           \a_mac_out[7]_cal1_u146_mac , \a_mac_out[7]_coefcal1_u63_mac ,
           \a_mac_out[7]_coefcal1_u64_mac , \a_mac_out[7]_coefcal1_u64_mac_0_ ,
           \a_mac_out[8]_cal1_u134_mac , \a_mac_out[8]_cal1_u135_mac , \a_mac_out[8]_cal1_u136_mac ,
           \a_mac_out[8]_cal1_u137_mac , \a_mac_out[8]_cal1_u138_mac , \a_mac_out[8]_cal1_u139_mac ,
           \a_mac_out[8]_cal1_u140_mac , \a_mac_out[8]_cal1_u141_mac , \a_mac_out[8]_cal1_u142_mac ,
           \a_mac_out[8]_cal1_u143_mac , \a_mac_out[8]_cal1_u144_mac , \a_mac_out[8]_cal1_u145_mac ,
           \a_mac_out[8]_cal1_u146_mac , \a_mac_out[8]_coefcal1_u63_mac ,
           \a_mac_out[8]_coefcal1_u64_mac , \a_mac_out[8]_coefcal1_u64_mac_0_ ,
           \a_mac_out[9]_cal1_u134_mac , \a_mac_out[9]_cal1_u135_mac , \a_mac_out[9]_cal1_u136_mac ,
           \a_mac_out[9]_cal1_u137_mac , \a_mac_out[9]_cal1_u138_mac , \a_mac_out[9]_cal1_u139_mac ,
           \a_mac_out[9]_cal1_u140_mac , \a_mac_out[9]_cal1_u141_mac , \a_mac_out[9]_cal1_u142_mac ,
           \a_mac_out[9]_cal1_u143_mac , \a_mac_out[9]_cal1_u144_mac , \a_mac_out[9]_cal1_u145_mac ,
           \a_mac_out[9]_cal1_u146_mac , \a_mac_out[9]_coefcal1_u63_mac ,
           \a_mac_out[9]_coefcal1_u64_mac , \a_mac_out[9]_coefcal1_u64_mac_0_ ,
           a_mac_out_cen_cal1_u134_mac, a_mac_out_cen_cal1_u135_mac, a_mac_out_cen_cal1_u136_mac,
           a_mac_out_cen_cal1_u137_mac, a_mac_out_cen_cal1_u138_mac, a_mac_out_cen_cal1_u139_mac,
           a_mac_out_cen_cal1_u140_mac, a_mac_out_cen_cal1_u141_mac, a_mac_out_cen_cal1_u142_mac,
           a_mac_out_cen_cal1_u143_mac, a_mac_out_cen_cal1_u144_mac, a_mac_out_cen_cal1_u145_mac,
           a_mac_out_cen_cal1_u146_mac, a_mac_out_cen_coefcal1_u63_mac, a_mac_out_cen_coefcal1_u64_mac,
           a_mac_out_cen_coefcal1_u64_mac_0_, a_out_sr_cal1_u134_mac, a_out_sr_cal1_u135_mac,
           a_out_sr_cal1_u136_mac, a_out_sr_cal1_u137_mac, a_out_sr_cal1_u138_mac,
           a_out_sr_cal1_u139_mac, a_out_sr_cal1_u140_mac, a_out_sr_cal1_u141_mac,
           a_out_sr_cal1_u142_mac, a_out_sr_cal1_u143_mac, a_out_sr_cal1_u144_mac,
           a_out_sr_cal1_u145_mac, a_out_sr_cal1_u146_mac, a_out_sr_coefcal1_u63_mac,
           a_out_sr_coefcal1_u64_mac, a_out_sr_coefcal1_u64_mac_0_, a_sload_cal1_u134_mac,
           a_sload_cal1_u135_mac, a_sload_cal1_u136_mac, a_sload_cal1_u137_mac,
           a_sload_cal1_u138_mac, a_sload_cal1_u139_mac, a_sload_cal1_u140_mac,
           a_sload_cal1_u141_mac, a_sload_cal1_u142_mac, a_sload_cal1_u143_mac,
           a_sload_cal1_u144_mac, a_sload_cal1_u145_mac, a_sload_cal1_u146_mac,
           a_sload_coefcal1_u63_mac, a_sload_coefcal1_u64_mac, a_sload_coefcal1_u64_mac_0_,
           b_acc_en_coefcal1_u64_mac, b_acc_en_coefcal1_u64_mac_0_, \b_dinx[0]_coefcal1_u64_mac ,
           \b_dinx[0]_coefcal1_u64_mac_0_ , \b_dinx[10]_coefcal1_u64_mac ,
           \b_dinx[10]_coefcal1_u64_mac_0_ , \b_dinx[11]_coefcal1_u64_mac ,
           \b_dinx[11]_coefcal1_u64_mac_0_ , \b_dinx[12]_coefcal1_u64_mac ,
           \b_dinx[12]_coefcal1_u64_mac_0_ , \b_dinx[13]_coefcal1_u64_mac ,
           \b_dinx[13]_coefcal1_u64_mac_0_ , \b_dinx[1]_coefcal1_u64_mac ,
           \b_dinx[1]_coefcal1_u64_mac_0_ , \b_dinx[2]_coefcal1_u64_mac ,
           \b_dinx[2]_coefcal1_u64_mac_0_ , \b_dinx[3]_coefcal1_u64_mac ,
           \b_dinx[3]_coefcal1_u64_mac_0_ , \b_dinx[4]_coefcal1_u64_mac ,
           \b_dinx[4]_coefcal1_u64_mac_0_ , \b_dinx[5]_coefcal1_u64_mac ,
           \b_dinx[5]_coefcal1_u64_mac_0_ , \b_dinx[6]_coefcal1_u64_mac ,
           \b_dinx[6]_coefcal1_u64_mac_0_ , \b_dinx[7]_coefcal1_u64_mac ,
           \b_dinx[7]_coefcal1_u64_mac_0_ , \b_dinx[8]_coefcal1_u64_mac ,
           \b_dinx[8]_coefcal1_u64_mac_0_ , \b_dinx[9]_coefcal1_u64_mac ,
           \b_dinx[9]_coefcal1_u64_mac_0_ , b_dinxy_cen_coefcal1_u64_mac,
           b_dinxy_cen_coefcal1_u64_mac_0_, \b_diny[0]_coefcal1_u64_mac ,
           \b_diny[0]_coefcal1_u64_mac_0_ , \b_diny[1]_coefcal1_u64_mac ,
           \b_diny[1]_coefcal1_u64_mac_0_ , \b_diny[2]_coefcal1_u64_mac ,
           \b_diny[2]_coefcal1_u64_mac_0_ , \b_diny[3]_coefcal1_u64_mac ,
           \b_diny[3]_coefcal1_u64_mac_0_ , \b_diny[4]_coefcal1_u64_mac ,
           \b_diny[4]_coefcal1_u64_mac_0_ , \b_diny[5]_coefcal1_u64_mac ,
           \b_diny[5]_coefcal1_u64_mac_0_ , \b_diny[6]_coefcal1_u64_mac ,
           \b_diny[6]_coefcal1_u64_mac_0_ , \b_diny[7]_coefcal1_u64_mac ,
           \b_diny[7]_coefcal1_u64_mac_0_ , \b_diny[8]_coefcal1_u64_mac ,
           \b_diny[8]_coefcal1_u64_mac_0_ , \b_diny[9]_coefcal1_u64_mac ,
           \b_diny[9]_coefcal1_u64_mac_0_ , b_dinz_cen_coefcal1_u64_mac, b_dinz_cen_coefcal1_u64_mac_0_,
           b_dinz_en_coefcal1_u64_mac, b_dinz_en_coefcal1_u64_mac_0_, b_in_sr_coefcal1_u64_mac,
           b_in_sr_coefcal1_u64_mac_0_, \b_mac_out[0]_coefcal1_u64_mac , \b_mac_out[1]_coefcal1_u64_mac ,
           \b_mac_out[2]_coefcal1_u64_mac , \b_mac_out[3]_coefcal1_u64_mac ,
           \b_mac_out[4]_coefcal1_u64_mac , b_mac_out_cen_coefcal1_u64_mac,
           b_mac_out_cen_coefcal1_u64_mac_0_, b_out_sr_coefcal1_u64_mac, b_out_sr_coefcal1_u64_mac_0_,
           b_sload_coefcal1_u64_mac, b_sload_coefcal1_u64_mac_0_, \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r1_clka_fifo1_ram_inst_0_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_0_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_1_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_2_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_3_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_0_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_1_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_2_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_3_u_emb18k_1, \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r1_rstna_fifo1_ram_inst_0_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_0_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_1_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_1_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_2_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_2_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_3_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_3_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_1, c1r2_clka_fifo1_ram_inst_0_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_0_u_emb18k_1, c1r2_clka_fifo1_ram_inst_1_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_1_u_emb18k_1, c1r2_clka_fifo1_ram_inst_2_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_2_u_emb18k_1, c1r2_clka_fifo1_ram_inst_3_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_3_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_0_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_0_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_1_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_1_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_2_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_2_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_3_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_3_u_emb18k_1, \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r2_rstna_fifo1_ram_inst_0_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_0_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_1_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_1_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_2_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_2_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_3_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_3_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_1, c1r3_clka_fifo1_ram_inst_0_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_0_u_emb18k_1, c1r3_clka_fifo1_ram_inst_1_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_1_u_emb18k_1, c1r3_clka_fifo1_ram_inst_2_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_2_u_emb18k_1, c1r3_clka_fifo1_ram_inst_3_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_3_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_0_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_0_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_1_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_1_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_2_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_2_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_3_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_3_u_emb18k_1, \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r3_rstna_fifo1_ram_inst_0_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_0_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_1_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_1_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_2_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_2_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_3_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_3_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_1, c1r4_clka_fifo1_ram_inst_0_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_0_u_emb18k_1, c1r4_clka_fifo1_ram_inst_1_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_1_u_emb18k_1, c1r4_clka_fifo1_ram_inst_2_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_2_u_emb18k_1, c1r4_clka_fifo1_ram_inst_3_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_3_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_0_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_0_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_1_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_1_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_2_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_2_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_3_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_3_u_emb18k_1, \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r4_rstna_fifo1_ram_inst_0_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_0_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_1_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_1_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_2_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_2_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_3_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_3_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_1, cea_fifo1_ram_inst_0_u_emb18k_0,
           cea_fifo1_ram_inst_0_u_emb18k_1, cea_fifo1_ram_inst_1_u_emb18k_0,
           cea_fifo1_ram_inst_1_u_emb18k_1, cea_fifo1_ram_inst_2_u_emb18k_0,
           cea_fifo1_ram_inst_2_u_emb18k_1, cea_fifo1_ram_inst_3_u_emb18k_0,
           cea_fifo1_ram_inst_3_u_emb18k_1, ceb_fifo1_ram_inst_0_u_emb18k_0,
           ceb_fifo1_ram_inst_0_u_emb18k_1, ceb_fifo1_ram_inst_1_u_emb18k_0,
           ceb_fifo1_ram_inst_1_u_emb18k_1, ceb_fifo1_ram_inst_2_u_emb18k_0,
           ceb_fifo1_ram_inst_2_u_emb18k_1, ceb_fifo1_ram_inst_3_u_emb18k_0,
           ceb_fifo1_ram_inst_3_u_emb18k_1, clka, clkb, dIn, dInEn, dOut,
           dOutEn, en, \haa[0]_fifo1_ram_inst_0_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_1_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_2_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_3_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_0_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_1_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_2_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_3_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_0_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_1_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_2_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_3_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_0_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_1_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_2_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_3_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3_u_emb18k_1 ,
           iHsyn, iVsyn, inXRes, inYRes, outXRes, outYRes, rst, u3634_OUT,
           u3662_O, u3662_O_4_, u3672_O, u4168_or2_41__I0, u4168_or2_41__I0_5_,
           u4168_or2_41__IN, u4510_I1, u6776_O, u6776_O_1_, u6776_O_2_, u6789_Y,
           u6796_O, u6810_D0, u6810_I0, u6810_I0_0_, u6810_I0_3_, u6810_IN,
           wea_fifo1_ram_inst_0_u_emb18k_0, wea_fifo1_ram_inst_0_u_emb18k_1,
           wea_fifo1_ram_inst_1_u_emb18k_0, wea_fifo1_ram_inst_1_u_emb18k_1,
           wea_fifo1_ram_inst_2_u_emb18k_0, wea_fifo1_ram_inst_2_u_emb18k_1,
           wea_fifo1_ram_inst_3_u_emb18k_0, wea_fifo1_ram_inst_3_u_emb18k_1,
           web_fifo1_ram_inst_0_u_emb18k_0, web_fifo1_ram_inst_0_u_emb18k_1,
           web_fifo1_ram_inst_1_u_emb18k_0, web_fifo1_ram_inst_1_u_emb18k_1,
           web_fifo1_ram_inst_2_u_emb18k_0, web_fifo1_ram_inst_2_u_emb18k_1,
           web_fifo1_ram_inst_3_u_emb18k_0, web_fifo1_ram_inst_3_u_emb18k_1,
           xBgn, xEnd, yBgn, yEnd );

    output HS, VS, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u135_mac, a_acc_en_cal1_u136_mac,
       a_acc_en_cal1_u137_mac, a_acc_en_cal1_u138_mac, a_acc_en_cal1_u139_mac,
       a_acc_en_cal1_u140_mac, a_acc_en_cal1_u141_mac, a_acc_en_cal1_u142_mac,
       a_acc_en_cal1_u143_mac, a_acc_en_cal1_u144_mac, a_acc_en_cal1_u145_mac,
       a_acc_en_cal1_u146_mac, a_acc_en_coefcal1_u63_mac, a_acc_en_coefcal1_u64_mac,
       a_acc_en_coefcal1_u64_mac_0_, \a_dinx[0]_cal1_u134_mac , \a_dinx[0]_cal1_u135_mac ,
       \a_dinx[0]_cal1_u136_mac , \a_dinx[0]_cal1_u137_mac , \a_dinx[0]_cal1_u138_mac ,
       \a_dinx[0]_cal1_u139_mac , \a_dinx[0]_cal1_u140_mac , \a_dinx[0]_cal1_u141_mac ,
       \a_dinx[0]_cal1_u142_mac , \a_dinx[0]_cal1_u143_mac , \a_dinx[0]_cal1_u144_mac ,
       \a_dinx[0]_cal1_u145_mac , \a_dinx[0]_cal1_u146_mac , \a_dinx[0]_coefcal1_u63_mac ,
       \a_dinx[0]_coefcal1_u64_mac , \a_dinx[0]_coefcal1_u64_mac_0_ , \a_dinx[10]_cal1_u134_mac ,
       \a_dinx[10]_cal1_u135_mac , \a_dinx[10]_cal1_u136_mac , \a_dinx[10]_cal1_u137_mac ,
       \a_dinx[10]_cal1_u138_mac , \a_dinx[10]_cal1_u139_mac , \a_dinx[10]_cal1_u140_mac ,
       \a_dinx[10]_cal1_u141_mac , \a_dinx[10]_cal1_u142_mac , \a_dinx[10]_cal1_u143_mac ,
       \a_dinx[10]_cal1_u144_mac , \a_dinx[10]_cal1_u145_mac , \a_dinx[10]_cal1_u146_mac ,
       \a_dinx[10]_coefcal1_u63_mac , \a_dinx[10]_coefcal1_u64_mac , \a_dinx[10]_coefcal1_u64_mac_0_ ,
       \a_dinx[11]_cal1_u134_mac , \a_dinx[11]_cal1_u135_mac , \a_dinx[11]_cal1_u136_mac ,
       \a_dinx[11]_cal1_u137_mac , \a_dinx[11]_cal1_u138_mac , \a_dinx[11]_cal1_u139_mac ,
       \a_dinx[11]_cal1_u140_mac , \a_dinx[11]_cal1_u141_mac , \a_dinx[11]_cal1_u142_mac ,
       \a_dinx[11]_cal1_u143_mac , \a_dinx[11]_cal1_u144_mac , \a_dinx[11]_cal1_u145_mac ,
       \a_dinx[11]_cal1_u146_mac , \a_dinx[11]_coefcal1_u63_mac , \a_dinx[11]_coefcal1_u64_mac ,
       \a_dinx[11]_coefcal1_u64_mac_0_ , \a_dinx[12]_cal1_u134_mac , \a_dinx[12]_cal1_u135_mac ,
       \a_dinx[12]_cal1_u136_mac , \a_dinx[12]_cal1_u137_mac , \a_dinx[12]_cal1_u138_mac ,
       \a_dinx[12]_cal1_u139_mac , \a_dinx[12]_cal1_u140_mac , \a_dinx[12]_cal1_u141_mac ,
       \a_dinx[12]_cal1_u142_mac , \a_dinx[12]_cal1_u143_mac , \a_dinx[12]_cal1_u144_mac ,
       \a_dinx[12]_cal1_u145_mac , \a_dinx[12]_cal1_u146_mac , \a_dinx[12]_coefcal1_u63_mac ,
       \a_dinx[12]_coefcal1_u64_mac , \a_dinx[12]_coefcal1_u64_mac_0_ , \a_dinx[13]_cal1_u134_mac ,
       \a_dinx[13]_cal1_u135_mac , \a_dinx[13]_cal1_u136_mac , \a_dinx[13]_cal1_u137_mac ,
       \a_dinx[13]_cal1_u138_mac , \a_dinx[13]_cal1_u139_mac , \a_dinx[13]_cal1_u140_mac ,
       \a_dinx[13]_cal1_u141_mac , \a_dinx[13]_cal1_u142_mac , \a_dinx[13]_cal1_u143_mac ,
       \a_dinx[13]_cal1_u144_mac , \a_dinx[13]_cal1_u145_mac , \a_dinx[13]_cal1_u146_mac ,
       \a_dinx[13]_coefcal1_u63_mac , \a_dinx[13]_coefcal1_u64_mac , \a_dinx[13]_coefcal1_u64_mac_0_ ,
       \a_dinx[1]_cal1_u134_mac , \a_dinx[1]_cal1_u135_mac , \a_dinx[1]_cal1_u136_mac ,
       \a_dinx[1]_cal1_u137_mac , \a_dinx[1]_cal1_u138_mac , \a_dinx[1]_cal1_u139_mac ,
       \a_dinx[1]_cal1_u140_mac , \a_dinx[1]_cal1_u141_mac , \a_dinx[1]_cal1_u142_mac ,
       \a_dinx[1]_cal1_u143_mac , \a_dinx[1]_cal1_u144_mac , \a_dinx[1]_cal1_u145_mac ,
       \a_dinx[1]_cal1_u146_mac , \a_dinx[1]_coefcal1_u63_mac , \a_dinx[1]_coefcal1_u64_mac ,
       \a_dinx[1]_coefcal1_u64_mac_0_ , \a_dinx[2]_cal1_u134_mac , \a_dinx[2]_cal1_u135_mac ,
       \a_dinx[2]_cal1_u136_mac , \a_dinx[2]_cal1_u137_mac , \a_dinx[2]_cal1_u138_mac ,
       \a_dinx[2]_cal1_u139_mac , \a_dinx[2]_cal1_u140_mac , \a_dinx[2]_cal1_u141_mac ,
       \a_dinx[2]_cal1_u142_mac , \a_dinx[2]_cal1_u143_mac , \a_dinx[2]_cal1_u144_mac ,
       \a_dinx[2]_cal1_u145_mac , \a_dinx[2]_cal1_u146_mac , \a_dinx[2]_coefcal1_u63_mac ,
       \a_dinx[2]_coefcal1_u64_mac , \a_dinx[2]_coefcal1_u64_mac_0_ , \a_dinx[3]_cal1_u134_mac ,
       \a_dinx[3]_cal1_u135_mac , \a_dinx[3]_cal1_u136_mac , \a_dinx[3]_cal1_u137_mac ,
       \a_dinx[3]_cal1_u138_mac , \a_dinx[3]_cal1_u139_mac , \a_dinx[3]_cal1_u140_mac ,
       \a_dinx[3]_cal1_u141_mac , \a_dinx[3]_cal1_u142_mac , \a_dinx[3]_cal1_u143_mac ,
       \a_dinx[3]_cal1_u144_mac , \a_dinx[3]_cal1_u145_mac , \a_dinx[3]_cal1_u146_mac ,
       \a_dinx[3]_coefcal1_u63_mac , \a_dinx[3]_coefcal1_u64_mac , \a_dinx[3]_coefcal1_u64_mac_0_ ,
       \a_dinx[4]_cal1_u134_mac , \a_dinx[4]_cal1_u135_mac , \a_dinx[4]_cal1_u136_mac ,
       \a_dinx[4]_cal1_u137_mac , \a_dinx[4]_cal1_u138_mac , \a_dinx[4]_cal1_u139_mac ,
       \a_dinx[4]_cal1_u140_mac , \a_dinx[4]_cal1_u141_mac , \a_dinx[4]_cal1_u142_mac ,
       \a_dinx[4]_cal1_u143_mac , \a_dinx[4]_cal1_u144_mac , \a_dinx[4]_cal1_u145_mac ,
       \a_dinx[4]_cal1_u146_mac , \a_dinx[4]_coefcal1_u63_mac , \a_dinx[4]_coefcal1_u64_mac ,
       \a_dinx[4]_coefcal1_u64_mac_0_ , \a_dinx[5]_cal1_u134_mac , \a_dinx[5]_cal1_u135_mac ,
       \a_dinx[5]_cal1_u136_mac , \a_dinx[5]_cal1_u137_mac , \a_dinx[5]_cal1_u138_mac ,
       \a_dinx[5]_cal1_u139_mac , \a_dinx[5]_cal1_u140_mac , \a_dinx[5]_cal1_u141_mac ,
       \a_dinx[5]_cal1_u142_mac , \a_dinx[5]_cal1_u143_mac , \a_dinx[5]_cal1_u144_mac ,
       \a_dinx[5]_cal1_u145_mac , \a_dinx[5]_cal1_u146_mac , \a_dinx[5]_coefcal1_u63_mac ,
       \a_dinx[5]_coefcal1_u64_mac , \a_dinx[5]_coefcal1_u64_mac_0_ , \a_dinx[6]_cal1_u134_mac ,
       \a_dinx[6]_cal1_u135_mac , \a_dinx[6]_cal1_u136_mac , \a_dinx[6]_cal1_u137_mac ,
       \a_dinx[6]_cal1_u138_mac , \a_dinx[6]_cal1_u139_mac , \a_dinx[6]_cal1_u140_mac ,
       \a_dinx[6]_cal1_u141_mac , \a_dinx[6]_cal1_u142_mac , \a_dinx[6]_cal1_u143_mac ,
       \a_dinx[6]_cal1_u144_mac , \a_dinx[6]_cal1_u145_mac , \a_dinx[6]_cal1_u146_mac ,
       \a_dinx[6]_coefcal1_u63_mac , \a_dinx[6]_coefcal1_u64_mac , \a_dinx[6]_coefcal1_u64_mac_0_ ,
       \a_dinx[7]_cal1_u134_mac , \a_dinx[7]_cal1_u135_mac , \a_dinx[7]_cal1_u136_mac ,
       \a_dinx[7]_cal1_u137_mac , \a_dinx[7]_cal1_u138_mac , \a_dinx[7]_cal1_u139_mac ,
       \a_dinx[7]_cal1_u140_mac , \a_dinx[7]_cal1_u141_mac , \a_dinx[7]_cal1_u142_mac ,
       \a_dinx[7]_cal1_u143_mac , \a_dinx[7]_cal1_u144_mac , \a_dinx[7]_cal1_u145_mac ,
       \a_dinx[7]_cal1_u146_mac , \a_dinx[7]_coefcal1_u63_mac , \a_dinx[7]_coefcal1_u64_mac ,
       \a_dinx[7]_coefcal1_u64_mac_0_ , \a_dinx[8]_cal1_u134_mac , \a_dinx[8]_cal1_u135_mac ,
       \a_dinx[8]_cal1_u136_mac , \a_dinx[8]_cal1_u137_mac , \a_dinx[8]_cal1_u138_mac ,
       \a_dinx[8]_cal1_u139_mac , \a_dinx[8]_cal1_u140_mac , \a_dinx[8]_cal1_u141_mac ,
       \a_dinx[8]_cal1_u142_mac , \a_dinx[8]_cal1_u143_mac , \a_dinx[8]_cal1_u144_mac ,
       \a_dinx[8]_cal1_u145_mac , \a_dinx[8]_cal1_u146_mac , \a_dinx[8]_coefcal1_u63_mac ,
       \a_dinx[8]_coefcal1_u64_mac , \a_dinx[8]_coefcal1_u64_mac_0_ , \a_dinx[9]_cal1_u134_mac ,
       \a_dinx[9]_cal1_u135_mac , \a_dinx[9]_cal1_u136_mac , \a_dinx[9]_cal1_u137_mac ,
       \a_dinx[9]_cal1_u138_mac , \a_dinx[9]_cal1_u139_mac , \a_dinx[9]_cal1_u140_mac ,
       \a_dinx[9]_cal1_u141_mac , \a_dinx[9]_cal1_u142_mac , \a_dinx[9]_cal1_u143_mac ,
       \a_dinx[9]_cal1_u144_mac , \a_dinx[9]_cal1_u145_mac , \a_dinx[9]_cal1_u146_mac ,
       \a_dinx[9]_coefcal1_u63_mac , \a_dinx[9]_coefcal1_u64_mac , \a_dinx[9]_coefcal1_u64_mac_0_ ,
       a_dinxy_cen_cal1_u134_mac, a_dinxy_cen_cal1_u135_mac, a_dinxy_cen_cal1_u136_mac,
       a_dinxy_cen_cal1_u137_mac, a_dinxy_cen_cal1_u138_mac, a_dinxy_cen_cal1_u139_mac,
       a_dinxy_cen_cal1_u140_mac, a_dinxy_cen_cal1_u141_mac, a_dinxy_cen_cal1_u142_mac,
       a_dinxy_cen_cal1_u143_mac, a_dinxy_cen_cal1_u144_mac, a_dinxy_cen_cal1_u145_mac,
       a_dinxy_cen_cal1_u146_mac, a_dinxy_cen_coefcal1_u63_mac, a_dinxy_cen_coefcal1_u64_mac,
       a_dinxy_cen_coefcal1_u64_mac_0_, \a_diny[0]_cal1_u134_mac , \a_diny[0]_cal1_u135_mac ,
       \a_diny[0]_cal1_u136_mac , \a_diny[0]_cal1_u137_mac , \a_diny[0]_cal1_u138_mac ,
       \a_diny[0]_cal1_u139_mac , \a_diny[0]_cal1_u140_mac , \a_diny[0]_cal1_u141_mac ,
       \a_diny[0]_cal1_u142_mac , \a_diny[0]_cal1_u143_mac , \a_diny[0]_cal1_u144_mac ,
       \a_diny[0]_cal1_u145_mac , \a_diny[0]_cal1_u146_mac , \a_diny[0]_coefcal1_u63_mac ,
       \a_diny[0]_coefcal1_u64_mac , \a_diny[0]_coefcal1_u64_mac_0_ , \a_diny[1]_cal1_u134_mac ,
       \a_diny[1]_cal1_u135_mac , \a_diny[1]_cal1_u136_mac , \a_diny[1]_cal1_u137_mac ,
       \a_diny[1]_cal1_u138_mac , \a_diny[1]_cal1_u139_mac , \a_diny[1]_cal1_u140_mac ,
       \a_diny[1]_cal1_u141_mac , \a_diny[1]_cal1_u142_mac , \a_diny[1]_cal1_u143_mac ,
       \a_diny[1]_cal1_u144_mac , \a_diny[1]_cal1_u145_mac , \a_diny[1]_cal1_u146_mac ,
       \a_diny[1]_coefcal1_u63_mac , \a_diny[1]_coefcal1_u64_mac , \a_diny[1]_coefcal1_u64_mac_0_ ,
       \a_diny[2]_cal1_u134_mac , \a_diny[2]_cal1_u135_mac , \a_diny[2]_cal1_u136_mac ,
       \a_diny[2]_cal1_u137_mac , \a_diny[2]_cal1_u138_mac , \a_diny[2]_cal1_u139_mac ,
       \a_diny[2]_cal1_u140_mac , \a_diny[2]_cal1_u141_mac , \a_diny[2]_cal1_u142_mac ,
       \a_diny[2]_cal1_u143_mac , \a_diny[2]_cal1_u144_mac , \a_diny[2]_cal1_u145_mac ,
       \a_diny[2]_cal1_u146_mac , \a_diny[2]_coefcal1_u63_mac , \a_diny[2]_coefcal1_u64_mac ,
       \a_diny[2]_coefcal1_u64_mac_0_ , \a_diny[3]_cal1_u134_mac , \a_diny[3]_cal1_u135_mac ,
       \a_diny[3]_cal1_u136_mac , \a_diny[3]_cal1_u137_mac , \a_diny[3]_cal1_u138_mac ,
       \a_diny[3]_cal1_u139_mac , \a_diny[3]_cal1_u140_mac , \a_diny[3]_cal1_u141_mac ,
       \a_diny[3]_cal1_u142_mac , \a_diny[3]_cal1_u143_mac , \a_diny[3]_cal1_u144_mac ,
       \a_diny[3]_cal1_u145_mac , \a_diny[3]_cal1_u146_mac , \a_diny[3]_coefcal1_u63_mac ,
       \a_diny[3]_coefcal1_u64_mac , \a_diny[3]_coefcal1_u64_mac_0_ , \a_diny[4]_cal1_u134_mac ,
       \a_diny[4]_cal1_u135_mac , \a_diny[4]_cal1_u136_mac , \a_diny[4]_cal1_u137_mac ,
       \a_diny[4]_cal1_u138_mac , \a_diny[4]_cal1_u139_mac , \a_diny[4]_cal1_u140_mac ,
       \a_diny[4]_cal1_u141_mac , \a_diny[4]_cal1_u142_mac , \a_diny[4]_cal1_u143_mac ,
       \a_diny[4]_cal1_u144_mac , \a_diny[4]_cal1_u145_mac , \a_diny[4]_cal1_u146_mac ,
       \a_diny[4]_coefcal1_u63_mac , \a_diny[4]_coefcal1_u64_mac , \a_diny[4]_coefcal1_u64_mac_0_ ,
       \a_diny[5]_cal1_u134_mac , \a_diny[5]_cal1_u135_mac , \a_diny[5]_cal1_u136_mac ,
       \a_diny[5]_cal1_u137_mac , \a_diny[5]_cal1_u138_mac , \a_diny[5]_cal1_u139_mac ,
       \a_diny[5]_cal1_u140_mac , \a_diny[5]_cal1_u141_mac , \a_diny[5]_cal1_u142_mac ,
       \a_diny[5]_cal1_u143_mac , \a_diny[5]_cal1_u144_mac , \a_diny[5]_cal1_u145_mac ,
       \a_diny[5]_cal1_u146_mac , \a_diny[5]_coefcal1_u63_mac , \a_diny[5]_coefcal1_u64_mac ,
       \a_diny[5]_coefcal1_u64_mac_0_ , \a_diny[6]_cal1_u134_mac , \a_diny[6]_cal1_u135_mac ,
       \a_diny[6]_cal1_u136_mac , \a_diny[6]_cal1_u137_mac , \a_diny[6]_cal1_u138_mac ,
       \a_diny[6]_cal1_u139_mac , \a_diny[6]_cal1_u140_mac , \a_diny[6]_cal1_u141_mac ,
       \a_diny[6]_cal1_u142_mac , \a_diny[6]_cal1_u143_mac , \a_diny[6]_cal1_u144_mac ,
       \a_diny[6]_cal1_u145_mac , \a_diny[6]_cal1_u146_mac , \a_diny[6]_coefcal1_u63_mac ,
       \a_diny[6]_coefcal1_u64_mac , \a_diny[6]_coefcal1_u64_mac_0_ , \a_diny[7]_cal1_u134_mac ,
       \a_diny[7]_cal1_u135_mac , \a_diny[7]_cal1_u136_mac , \a_diny[7]_cal1_u137_mac ,
       \a_diny[7]_cal1_u138_mac , \a_diny[7]_cal1_u139_mac , \a_diny[7]_cal1_u140_mac ,
       \a_diny[7]_cal1_u141_mac , \a_diny[7]_cal1_u142_mac , \a_diny[7]_cal1_u143_mac ,
       \a_diny[7]_cal1_u144_mac , \a_diny[7]_cal1_u145_mac , \a_diny[7]_cal1_u146_mac ,
       \a_diny[7]_coefcal1_u63_mac , \a_diny[7]_coefcal1_u64_mac , \a_diny[7]_coefcal1_u64_mac_0_ ,
       \a_diny[8]_cal1_u134_mac , \a_diny[8]_cal1_u135_mac , \a_diny[8]_cal1_u136_mac ,
       \a_diny[8]_cal1_u137_mac , \a_diny[8]_cal1_u138_mac , \a_diny[8]_cal1_u139_mac ,
       \a_diny[8]_cal1_u140_mac , \a_diny[8]_cal1_u141_mac , \a_diny[8]_cal1_u142_mac ,
       \a_diny[8]_cal1_u143_mac , \a_diny[8]_cal1_u144_mac , \a_diny[8]_cal1_u145_mac ,
       \a_diny[8]_cal1_u146_mac , \a_diny[8]_coefcal1_u63_mac , \a_diny[8]_coefcal1_u64_mac ,
       \a_diny[8]_coefcal1_u64_mac_0_ , \a_diny[9]_cal1_u134_mac , \a_diny[9]_cal1_u135_mac ,
       \a_diny[9]_cal1_u136_mac , \a_diny[9]_cal1_u137_mac , \a_diny[9]_cal1_u138_mac ,
       \a_diny[9]_cal1_u139_mac , \a_diny[9]_cal1_u140_mac , \a_diny[9]_cal1_u141_mac ,
       \a_diny[9]_cal1_u142_mac , \a_diny[9]_cal1_u143_mac , \a_diny[9]_cal1_u144_mac ,
       \a_diny[9]_cal1_u145_mac , \a_diny[9]_cal1_u146_mac , \a_diny[9]_coefcal1_u63_mac ,
       \a_diny[9]_coefcal1_u64_mac , \a_diny[9]_coefcal1_u64_mac_0_ , a_dinz_cen_cal1_u134_mac,
       a_dinz_cen_cal1_u135_mac, a_dinz_cen_cal1_u136_mac, a_dinz_cen_cal1_u137_mac,
       a_dinz_cen_cal1_u138_mac, a_dinz_cen_cal1_u139_mac, a_dinz_cen_cal1_u140_mac,
       a_dinz_cen_cal1_u141_mac, a_dinz_cen_cal1_u142_mac, a_dinz_cen_cal1_u143_mac,
       a_dinz_cen_cal1_u144_mac, a_dinz_cen_cal1_u145_mac, a_dinz_cen_cal1_u146_mac,
       a_dinz_cen_coefcal1_u63_mac, a_dinz_cen_coefcal1_u64_mac, a_dinz_cen_coefcal1_u64_mac_0_,
       a_dinz_en_cal1_u134_mac, a_dinz_en_cal1_u135_mac, a_dinz_en_cal1_u136_mac,
       a_dinz_en_cal1_u137_mac, a_dinz_en_cal1_u138_mac, a_dinz_en_cal1_u139_mac,
       a_dinz_en_cal1_u140_mac, a_dinz_en_cal1_u141_mac, a_dinz_en_cal1_u142_mac,
       a_dinz_en_cal1_u143_mac, a_dinz_en_cal1_u144_mac, a_dinz_en_cal1_u145_mac,
       a_dinz_en_cal1_u146_mac, a_dinz_en_coefcal1_u63_mac, a_dinz_en_coefcal1_u64_mac,
       a_dinz_en_coefcal1_u64_mac_0_, a_in_sr_cal1_u134_mac, a_in_sr_cal1_u135_mac,
       a_in_sr_cal1_u136_mac, a_in_sr_cal1_u137_mac, a_in_sr_cal1_u138_mac, a_in_sr_cal1_u139_mac,
       a_in_sr_cal1_u140_mac, a_in_sr_cal1_u141_mac, a_in_sr_cal1_u142_mac, a_in_sr_cal1_u143_mac,
       a_in_sr_cal1_u144_mac, a_in_sr_cal1_u145_mac, a_in_sr_cal1_u146_mac, a_in_sr_coefcal1_u63_mac,
       a_in_sr_coefcal1_u64_mac, a_in_sr_coefcal1_u64_mac_0_;
    input  \a_mac_out[0]_coefcal1_u63_mac , \a_mac_out[0]_coefcal1_u64_mac ,
       \a_mac_out[0]_coefcal1_u64_mac_0_ , \a_mac_out[10]_cal1_u134_mac , \a_mac_out[10]_cal1_u135_mac ,
       \a_mac_out[10]_cal1_u136_mac , \a_mac_out[10]_cal1_u137_mac , \a_mac_out[10]_cal1_u138_mac ,
       \a_mac_out[10]_cal1_u139_mac , \a_mac_out[10]_cal1_u140_mac , \a_mac_out[10]_cal1_u141_mac ,
       \a_mac_out[10]_cal1_u142_mac , \a_mac_out[10]_cal1_u143_mac , \a_mac_out[10]_cal1_u144_mac ,
       \a_mac_out[10]_cal1_u145_mac , \a_mac_out[10]_cal1_u146_mac , \a_mac_out[10]_coefcal1_u63_mac ,
       \a_mac_out[10]_coefcal1_u64_mac , \a_mac_out[10]_coefcal1_u64_mac_0_ ,
       \a_mac_out[11]_cal1_u134_mac , \a_mac_out[11]_cal1_u139_mac , \a_mac_out[11]_cal1_u140_mac ,
       \a_mac_out[11]_cal1_u141_mac , \a_mac_out[11]_cal1_u142_mac , \a_mac_out[11]_coefcal1_u63_mac ,
       \a_mac_out[11]_coefcal1_u64_mac , \a_mac_out[11]_coefcal1_u64_mac_0_ ,
       \a_mac_out[12]_coefcal1_u63_mac , \a_mac_out[12]_coefcal1_u64_mac , \a_mac_out[12]_coefcal1_u64_mac_0_ ,
       \a_mac_out[13]_coefcal1_u63_mac , \a_mac_out[13]_coefcal1_u64_mac , \a_mac_out[14]_coefcal1_u63_mac ,
       \a_mac_out[14]_coefcal1_u64_mac , \a_mac_out[15]_coefcal1_u63_mac , \a_mac_out[15]_coefcal1_u64_mac ,
       \a_mac_out[16]_coefcal1_u63_mac , \a_mac_out[16]_coefcal1_u64_mac , \a_mac_out[17]_coefcal1_u63_mac ,
       \a_mac_out[17]_coefcal1_u64_mac , \a_mac_out[18]_coefcal1_u63_mac , \a_mac_out[18]_coefcal1_u64_mac ,
       \a_mac_out[19]_coefcal1_u63_mac , \a_mac_out[19]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u63_mac ,
       \a_mac_out[1]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u64_mac_0_ , \a_mac_out[20]_coefcal1_u64_mac ,
       \a_mac_out[21]_coefcal1_u64_mac , \a_mac_out[22]_coefcal1_u64_mac , \a_mac_out[23]_coefcal1_u64_mac ,
       \a_mac_out[2]_coefcal1_u63_mac , \a_mac_out[2]_coefcal1_u64_mac , \a_mac_out[2]_coefcal1_u64_mac_0_ ,
       \a_mac_out[3]_coefcal1_u63_mac , \a_mac_out[3]_coefcal1_u64_mac , \a_mac_out[3]_coefcal1_u64_mac_0_ ,
       \a_mac_out[4]_coefcal1_u63_mac , \a_mac_out[4]_coefcal1_u64_mac , \a_mac_out[4]_coefcal1_u64_mac_0_ ,
       \a_mac_out[5]_coefcal1_u63_mac , \a_mac_out[5]_coefcal1_u64_mac , \a_mac_out[5]_coefcal1_u64_mac_0_ ,
       \a_mac_out[6]_cal1_u134_mac , \a_mac_out[6]_cal1_u135_mac , \a_mac_out[6]_cal1_u136_mac ,
       \a_mac_out[6]_cal1_u137_mac , \a_mac_out[6]_cal1_u138_mac , \a_mac_out[6]_cal1_u139_mac ,
       \a_mac_out[6]_cal1_u140_mac , \a_mac_out[6]_cal1_u141_mac , \a_mac_out[6]_cal1_u142_mac ,
       \a_mac_out[6]_cal1_u143_mac , \a_mac_out[6]_cal1_u144_mac , \a_mac_out[6]_cal1_u145_mac ,
       \a_mac_out[6]_cal1_u146_mac , \a_mac_out[6]_coefcal1_u63_mac , \a_mac_out[6]_coefcal1_u64_mac ,
       \a_mac_out[6]_coefcal1_u64_mac_0_ , \a_mac_out[7]_cal1_u134_mac , \a_mac_out[7]_cal1_u135_mac ,
       \a_mac_out[7]_cal1_u136_mac , \a_mac_out[7]_cal1_u137_mac , \a_mac_out[7]_cal1_u138_mac ,
       \a_mac_out[7]_cal1_u139_mac , \a_mac_out[7]_cal1_u140_mac , \a_mac_out[7]_cal1_u141_mac ,
       \a_mac_out[7]_cal1_u142_mac , \a_mac_out[7]_cal1_u143_mac , \a_mac_out[7]_cal1_u144_mac ,
       \a_mac_out[7]_cal1_u145_mac , \a_mac_out[7]_cal1_u146_mac , \a_mac_out[7]_coefcal1_u63_mac ,
       \a_mac_out[7]_coefcal1_u64_mac , \a_mac_out[7]_coefcal1_u64_mac_0_ , \a_mac_out[8]_cal1_u134_mac ,
       \a_mac_out[8]_cal1_u135_mac , \a_mac_out[8]_cal1_u136_mac , \a_mac_out[8]_cal1_u137_mac ,
       \a_mac_out[8]_cal1_u138_mac , \a_mac_out[8]_cal1_u139_mac , \a_mac_out[8]_cal1_u140_mac ,
       \a_mac_out[8]_cal1_u141_mac , \a_mac_out[8]_cal1_u142_mac , \a_mac_out[8]_cal1_u143_mac ,
       \a_mac_out[8]_cal1_u144_mac , \a_mac_out[8]_cal1_u145_mac , \a_mac_out[8]_cal1_u146_mac ,
       \a_mac_out[8]_coefcal1_u63_mac , \a_mac_out[8]_coefcal1_u64_mac , \a_mac_out[8]_coefcal1_u64_mac_0_ ,
       \a_mac_out[9]_cal1_u134_mac , \a_mac_out[9]_cal1_u135_mac , \a_mac_out[9]_cal1_u136_mac ,
       \a_mac_out[9]_cal1_u137_mac , \a_mac_out[9]_cal1_u138_mac , \a_mac_out[9]_cal1_u139_mac ,
       \a_mac_out[9]_cal1_u140_mac , \a_mac_out[9]_cal1_u141_mac , \a_mac_out[9]_cal1_u142_mac ,
       \a_mac_out[9]_cal1_u143_mac , \a_mac_out[9]_cal1_u144_mac , \a_mac_out[9]_cal1_u145_mac ,
       \a_mac_out[9]_cal1_u146_mac , \a_mac_out[9]_coefcal1_u63_mac , \a_mac_out[9]_coefcal1_u64_mac ,
       \a_mac_out[9]_coefcal1_u64_mac_0_ ;
    output a_mac_out_cen_cal1_u134_mac, a_mac_out_cen_cal1_u135_mac, a_mac_out_cen_cal1_u136_mac,
       a_mac_out_cen_cal1_u137_mac, a_mac_out_cen_cal1_u138_mac, a_mac_out_cen_cal1_u139_mac,
       a_mac_out_cen_cal1_u140_mac, a_mac_out_cen_cal1_u141_mac, a_mac_out_cen_cal1_u142_mac,
       a_mac_out_cen_cal1_u143_mac, a_mac_out_cen_cal1_u144_mac, a_mac_out_cen_cal1_u145_mac,
       a_mac_out_cen_cal1_u146_mac, a_mac_out_cen_coefcal1_u63_mac, a_mac_out_cen_coefcal1_u64_mac,
       a_mac_out_cen_coefcal1_u64_mac_0_, a_out_sr_cal1_u134_mac, a_out_sr_cal1_u135_mac,
       a_out_sr_cal1_u136_mac, a_out_sr_cal1_u137_mac, a_out_sr_cal1_u138_mac,
       a_out_sr_cal1_u139_mac, a_out_sr_cal1_u140_mac, a_out_sr_cal1_u141_mac,
       a_out_sr_cal1_u142_mac, a_out_sr_cal1_u143_mac, a_out_sr_cal1_u144_mac,
       a_out_sr_cal1_u145_mac, a_out_sr_cal1_u146_mac, a_out_sr_coefcal1_u63_mac,
       a_out_sr_coefcal1_u64_mac, a_out_sr_coefcal1_u64_mac_0_, a_sload_cal1_u134_mac,
       a_sload_cal1_u135_mac, a_sload_cal1_u136_mac, a_sload_cal1_u137_mac, a_sload_cal1_u138_mac,
       a_sload_cal1_u139_mac, a_sload_cal1_u140_mac, a_sload_cal1_u141_mac, a_sload_cal1_u142_mac,
       a_sload_cal1_u143_mac, a_sload_cal1_u144_mac, a_sload_cal1_u145_mac, a_sload_cal1_u146_mac,
       a_sload_coefcal1_u63_mac, a_sload_coefcal1_u64_mac, a_sload_coefcal1_u64_mac_0_,
       b_acc_en_coefcal1_u64_mac, b_acc_en_coefcal1_u64_mac_0_, \b_dinx[0]_coefcal1_u64_mac ,
       \b_dinx[0]_coefcal1_u64_mac_0_ , \b_dinx[10]_coefcal1_u64_mac , \b_dinx[10]_coefcal1_u64_mac_0_ ,
       \b_dinx[11]_coefcal1_u64_mac , \b_dinx[11]_coefcal1_u64_mac_0_ , \b_dinx[12]_coefcal1_u64_mac ,
       \b_dinx[12]_coefcal1_u64_mac_0_ , \b_dinx[13]_coefcal1_u64_mac , \b_dinx[13]_coefcal1_u64_mac_0_ ,
       \b_dinx[1]_coefcal1_u64_mac , \b_dinx[1]_coefcal1_u64_mac_0_ , \b_dinx[2]_coefcal1_u64_mac ,
       \b_dinx[2]_coefcal1_u64_mac_0_ , \b_dinx[3]_coefcal1_u64_mac , \b_dinx[3]_coefcal1_u64_mac_0_ ,
       \b_dinx[4]_coefcal1_u64_mac , \b_dinx[4]_coefcal1_u64_mac_0_ , \b_dinx[5]_coefcal1_u64_mac ,
       \b_dinx[5]_coefcal1_u64_mac_0_ , \b_dinx[6]_coefcal1_u64_mac , \b_dinx[6]_coefcal1_u64_mac_0_ ,
       \b_dinx[7]_coefcal1_u64_mac , \b_dinx[7]_coefcal1_u64_mac_0_ , \b_dinx[8]_coefcal1_u64_mac ,
       \b_dinx[8]_coefcal1_u64_mac_0_ , \b_dinx[9]_coefcal1_u64_mac , \b_dinx[9]_coefcal1_u64_mac_0_ ,
       b_dinxy_cen_coefcal1_u64_mac, b_dinxy_cen_coefcal1_u64_mac_0_, \b_diny[0]_coefcal1_u64_mac ,
       \b_diny[0]_coefcal1_u64_mac_0_ , \b_diny[1]_coefcal1_u64_mac , \b_diny[1]_coefcal1_u64_mac_0_ ,
       \b_diny[2]_coefcal1_u64_mac , \b_diny[2]_coefcal1_u64_mac_0_ , \b_diny[3]_coefcal1_u64_mac ,
       \b_diny[3]_coefcal1_u64_mac_0_ , \b_diny[4]_coefcal1_u64_mac , \b_diny[4]_coefcal1_u64_mac_0_ ,
       \b_diny[5]_coefcal1_u64_mac , \b_diny[5]_coefcal1_u64_mac_0_ , \b_diny[6]_coefcal1_u64_mac ,
       \b_diny[6]_coefcal1_u64_mac_0_ , \b_diny[7]_coefcal1_u64_mac , \b_diny[7]_coefcal1_u64_mac_0_ ,
       \b_diny[8]_coefcal1_u64_mac , \b_diny[8]_coefcal1_u64_mac_0_ , \b_diny[9]_coefcal1_u64_mac ,
       \b_diny[9]_coefcal1_u64_mac_0_ , b_dinz_cen_coefcal1_u64_mac, b_dinz_cen_coefcal1_u64_mac_0_,
       b_dinz_en_coefcal1_u64_mac, b_dinz_en_coefcal1_u64_mac_0_, b_in_sr_coefcal1_u64_mac,
       b_in_sr_coefcal1_u64_mac_0_;
    input  \b_mac_out[0]_coefcal1_u64_mac , \b_mac_out[1]_coefcal1_u64_mac ,
       \b_mac_out[2]_coefcal1_u64_mac , \b_mac_out[3]_coefcal1_u64_mac , \b_mac_out[4]_coefcal1_u64_mac ;
    output b_mac_out_cen_coefcal1_u64_mac, b_mac_out_cen_coefcal1_u64_mac_0_,
       b_out_sr_coefcal1_u64_mac, b_out_sr_coefcal1_u64_mac_0_, b_sload_coefcal1_u64_mac,
       b_sload_coefcal1_u64_mac_0_, \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_1 , c1r1_clka_fifo1_ram_inst_0_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_0_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_1_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_2_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_3_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_0_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_1_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_2_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_3_u_emb18k_1, \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    input  \c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    output c1r1_rstna_fifo1_ram_inst_0_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_0_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_1_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_1_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_2_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_2_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_3_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_3_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_0_u_emb18k_0, c1r2_clka_fifo1_ram_inst_0_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_1_u_emb18k_0, c1r2_clka_fifo1_ram_inst_1_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_2_u_emb18k_0, c1r2_clka_fifo1_ram_inst_2_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_3_u_emb18k_0, c1r2_clka_fifo1_ram_inst_3_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_0_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_0_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_1_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_1_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_2_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_2_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_3_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_3_u_emb18k_1,
       \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    input  \c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    output c1r2_rstna_fifo1_ram_inst_0_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_0_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_1_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_1_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_2_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_2_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_3_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_3_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_0_u_emb18k_0, c1r3_clka_fifo1_ram_inst_0_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_1_u_emb18k_0, c1r3_clka_fifo1_ram_inst_1_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_2_u_emb18k_0, c1r3_clka_fifo1_ram_inst_2_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_3_u_emb18k_0, c1r3_clka_fifo1_ram_inst_3_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_0_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_0_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_1_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_1_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_2_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_2_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_3_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_3_u_emb18k_1,
       \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    input  \c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    output c1r3_rstna_fifo1_ram_inst_0_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_0_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_1_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_1_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_2_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_2_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_3_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_3_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_0_u_emb18k_0, c1r4_clka_fifo1_ram_inst_0_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_1_u_emb18k_0, c1r4_clka_fifo1_ram_inst_1_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_2_u_emb18k_0, c1r4_clka_fifo1_ram_inst_2_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_3_u_emb18k_0, c1r4_clka_fifo1_ram_inst_3_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_0_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_0_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_1_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_1_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_2_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_2_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_3_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_3_u_emb18k_1,
       \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    input  \c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_1 ,
       \c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_1 ,
       \c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_1 ,
       \c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_1 ;
    output c1r4_rstna_fifo1_ram_inst_0_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_0_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_1_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_1_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_2_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_2_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_3_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_3_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_1,
       cea_fifo1_ram_inst_0_u_emb18k_0, cea_fifo1_ram_inst_0_u_emb18k_1, cea_fifo1_ram_inst_1_u_emb18k_0,
       cea_fifo1_ram_inst_1_u_emb18k_1, cea_fifo1_ram_inst_2_u_emb18k_0, cea_fifo1_ram_inst_2_u_emb18k_1,
       cea_fifo1_ram_inst_3_u_emb18k_0, cea_fifo1_ram_inst_3_u_emb18k_1, ceb_fifo1_ram_inst_0_u_emb18k_0,
       ceb_fifo1_ram_inst_0_u_emb18k_1, ceb_fifo1_ram_inst_1_u_emb18k_0, ceb_fifo1_ram_inst_1_u_emb18k_1,
       ceb_fifo1_ram_inst_2_u_emb18k_0, ceb_fifo1_ram_inst_2_u_emb18k_1, ceb_fifo1_ram_inst_3_u_emb18k_0,
       ceb_fifo1_ram_inst_3_u_emb18k_1;
    input  clka, clkb;
    input  [15:0] dIn;
    input  dInEn;
    output [15:0] dOut;
    output dOutEn;
    input  en;
    output \haa[0]_fifo1_ram_inst_0_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_1_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_2_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_3_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_0_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_1_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_2_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_3_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_0_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_1_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_2_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_3_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_0_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_1_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_2_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_3_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3_u_emb18k_1 ;
    input  iHsyn, iVsyn;
    input  [10:0] inXRes;
    input  [10:0] inYRes;
    input  [11:0] outXRes;
    input  [11:0] outYRes;
    input  rst;
    output u3634_OUT, u3662_O, u3662_O_4_, u3672_O;
    input  u4168_or2_41__I0, u4168_or2_41__I0_5_, u4168_or2_41__IN, u4510_I1;
    output u6776_O, u6776_O_1_, u6776_O_2_, u6789_Y, u6796_O;
    input  u6810_D0, u6810_I0, u6810_I0_0_, u6810_I0_3_, u6810_IN;
    output wea_fifo1_ram_inst_0_u_emb18k_0, wea_fifo1_ram_inst_0_u_emb18k_1,
       wea_fifo1_ram_inst_1_u_emb18k_0, wea_fifo1_ram_inst_1_u_emb18k_1, wea_fifo1_ram_inst_2_u_emb18k_0,
       wea_fifo1_ram_inst_2_u_emb18k_1, wea_fifo1_ram_inst_3_u_emb18k_0, wea_fifo1_ram_inst_3_u_emb18k_1,
       web_fifo1_ram_inst_0_u_emb18k_0, web_fifo1_ram_inst_0_u_emb18k_1, web_fifo1_ram_inst_1_u_emb18k_0,
       web_fifo1_ram_inst_1_u_emb18k_1, web_fifo1_ram_inst_2_u_emb18k_0, web_fifo1_ram_inst_2_u_emb18k_1,
       web_fifo1_ram_inst_3_u_emb18k_0, web_fifo1_ram_inst_3_u_emb18k_1;
    input  [10:0] xBgn;
    input  [10:0] xEnd;
    input  [10:0] yBgn;
    input  [10:0] yEnd;
    wire   HS_1863_net, \cal1_VSNormal__reg|Q_net , \cal1_enforceJmp__reg|Q_net ,
       \cal1_jmp1Normal__reg|Q_net , \cal1_jmp2Normal__reg|Q_net , \cal1_ramRdAddr__reg[0]|Q_net ,
       \cal1_ramRdAddr__reg[10]|Q_net , \cal1_ramRdAddr__reg[1]|Q_net , \cal1_ramRdAddr__reg[2]|Q_net ,
       \cal1_ramRdAddr__reg[3]|Q_net , \cal1_ramRdAddr__reg[4]|Q_net , \cal1_ramRdAddr__reg[5]|Q_net ,
       \cal1_ramRdAddr__reg[6]|Q_net , \cal1_ramRdAddr__reg[7]|Q_net , \cal1_ramRdAddr__reg[8]|Q_net ,
       \cal1_ramRdAddr__reg[9]|Q_net , \cal1_u127_XORCI_0|SUM_net , \cal1_u127_XORCI_10|SUM_net ,
       \cal1_u127_XORCI_11|SUM_net , \cal1_u127_XORCI_12|SUM_net , \cal1_u127_XORCI_13|SUM_net ,
       \cal1_u127_XORCI_14|SUM_net , \cal1_u127_XORCI_15|SUM_net , \cal1_u127_XORCI_16|SUM_net ,
       \cal1_u127_XORCI_1|SUM_net , \cal1_u127_XORCI_2|SUM_net , \cal1_u127_XORCI_3|SUM_net ,
       \cal1_u127_XORCI_4|SUM_net , \cal1_u127_XORCI_5|SUM_net , \cal1_u127_XORCI_6|SUM_net ,
       \cal1_u127_XORCI_7|SUM_net , \cal1_u127_XORCI_8|SUM_net , \cal1_u127_XORCI_9|SUM_net ,
       \cal1_u128_XORCI_0|SUM_net , \cal1_u128_XORCI_10|SUM_net , \cal1_u128_XORCI_11|SUM_net ,
       \cal1_u128_XORCI_12|SUM_net , \cal1_u128_XORCI_13|SUM_net , \cal1_u128_XORCI_14|SUM_net ,
       \cal1_u128_XORCI_15|SUM_net , \cal1_u128_XORCI_16|SUM_net , \cal1_u128_XORCI_1|SUM_net ,
       \cal1_u128_XORCI_2|SUM_net , \cal1_u128_XORCI_3|SUM_net , \cal1_u128_XORCI_4|SUM_net ,
       \cal1_u128_XORCI_5|SUM_net , \cal1_u128_XORCI_6|SUM_net , \cal1_u128_XORCI_7|SUM_net ,
       \cal1_u128_XORCI_8|SUM_net , \cal1_u128_XORCI_9|SUM_net , \cal1_u129_XORCI_0|SUM_net ,
       \cal1_u129_XORCI_10|SUM_net , \cal1_u129_XORCI_1|SUM_net , \cal1_u129_XORCI_2|SUM_net ,
       \cal1_u129_XORCI_3|SUM_net , \cal1_u129_XORCI_4|SUM_net , \cal1_u129_XORCI_5|SUM_net ,
       \cal1_u129_XORCI_6|SUM_net , \cal1_u129_XORCI_7|SUM_net , \cal1_u129_XORCI_8|SUM_net ,
       \cal1_u129_XORCI_9|SUM_net , \cal1_u130_XORCI_0|SUM_net , \cal1_u130_XORCI_10|SUM_net ,
       \cal1_u130_XORCI_1|SUM_net , \cal1_u130_XORCI_2|SUM_net , \cal1_u130_XORCI_3|SUM_net ,
       \cal1_u130_XORCI_4|SUM_net , \cal1_u130_XORCI_5|SUM_net , \cal1_u130_XORCI_6|SUM_net ,
       \cal1_u130_XORCI_7|SUM_net , \cal1_u130_XORCI_8|SUM_net , \cal1_u130_XORCI_9|SUM_net ,
       \cal1_u131_XORCI_0|SUM_net , \cal1_u131_XORCI_10|SUM_net , \cal1_u131_XORCI_1|SUM_net ,
       \cal1_u131_XORCI_2|SUM_net , \cal1_u131_XORCI_3|SUM_net , \cal1_u131_XORCI_4|SUM_net ,
       \cal1_u131_XORCI_5|SUM_net , \cal1_u131_XORCI_6|SUM_net , \cal1_u131_XORCI_7|SUM_net ,
       \cal1_u131_XORCI_8|SUM_net , \cal1_u131_XORCI_9|SUM_net , \cal1_u132_XORCI_0|SUM_net ,
       \cal1_u132_XORCI_10|SUM_net , \cal1_u132_XORCI_1|SUM_net , \cal1_u132_XORCI_2|SUM_net ,
       \cal1_u132_XORCI_3|SUM_net , \cal1_u132_XORCI_4|SUM_net , \cal1_u132_XORCI_5|SUM_net ,
       \cal1_u132_XORCI_6|SUM_net , \cal1_u132_XORCI_7|SUM_net , \cal1_u132_XORCI_8|SUM_net ,
       \cal1_u132_XORCI_9|SUM_net , \cal1_u133_XORCI_0|SUM_net , \cal1_u133_XORCI_1|SUM_net ,
       \cal1_u133_XORCI_2|SUM_net , \cal1_u133_XORCI_3|SUM_net , \cal1_u133_XORCI_4|SUM_net ,
       \cal1_u133_XORCI_5|SUM_net , \cal1_u133_XORCI_6|SUM_net , \cal1_u54_XORCI_0|SUM_net ,
       \cal1_u54_XORCI_1|SUM_net , \cal1_u54_XORCI_2|SUM_net , \cal1_u54_XORCI_3|SUM_net ,
       \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_5|SUM_net , \cal1_u54_XORCI_6|SUM_net ,
       \cal1_u55_XORCI_0|SUM_net , \cal1_u55_XORCI_1|SUM_net , \cal1_u55_XORCI_2|SUM_net ,
       \cal1_u55_XORCI_3|SUM_net , \cal1_u55_XORCI_4|SUM_net , \cal1_u55_XORCI_5|SUM_net ,
       \cal1_u55_XORCI_6|SUM_net , \cal1_u57_XORCI_11|SUM_net , \cal1_u59_XORCI_11|SUM_net ,
       \cal1_u61_XORCI_11|SUM_net , \cal1_u63_XORCI_11|SUM_net , \cal1_uPreF__reg[0]|Q_net ,
       \cal1_uPreF__reg[1]|Q_net , \cal1_uPreF__reg[2]|Q_net , \cal1_uPreF__reg[3]|Q_net ,
       \cal1_uPreF__reg[4]|Q_net , \cal1_uPreF__reg[5]|Q_net , \cal1_u__reg[0]|Q_net ,
       \cal1_u__reg[10]|Q_net , \cal1_u__reg[11]|Q_net , \cal1_u__reg[12]|Q_net ,
       \cal1_u__reg[13]|Q_net , \cal1_u__reg[14]|Q_net , \cal1_u__reg[15]|Q_net ,
       \cal1_u__reg[16]|Q_net , \cal1_u__reg[1]|Q_net , \cal1_u__reg[2]|Q_net ,
       \cal1_u__reg[3]|Q_net , \cal1_u__reg[4]|Q_net , \cal1_u__reg[5]|Q_net ,
       \cal1_u__reg[6]|Q_net , \cal1_u__reg[7]|Q_net , \cal1_u__reg[8]|Q_net ,
       \cal1_u__reg[9]|Q_net , \cal1_v__reg[0]|Q_net , \cal1_v__reg[10]|Q_net ,
       \cal1_v__reg[11]|Q_net , \cal1_v__reg[12]|Q_net , \cal1_v__reg[13]|Q_net ,
       \cal1_v__reg[14]|Q_net , \cal1_v__reg[15]|Q_net , \cal1_v__reg[16]|Q_net ,
       \cal1_v__reg[1]|Q_net , \cal1_v__reg[2]|Q_net , \cal1_v__reg[3]|Q_net ,
       \cal1_v__reg[4]|Q_net , \cal1_v__reg[5]|Q_net , \cal1_v__reg[6]|Q_net ,
       \cal1_v__reg[7]|Q_net , \cal1_v__reg[8]|Q_net , \cal1_v__reg[9]|Q_net ,
       \cal1_xAddress__reg[0]|Q_net , \cal1_xAddress__reg[10]|Q_net , \cal1_xAddress__reg[1]|Q_net ,
       \cal1_xAddress__reg[2]|Q_net , \cal1_xAddress__reg[3]|Q_net , \cal1_xAddress__reg[4]|Q_net ,
       \cal1_xAddress__reg[5]|Q_net , \cal1_xAddress__reg[6]|Q_net , \cal1_xAddress__reg[7]|Q_net ,
       \cal1_xAddress__reg[8]|Q_net , \cal1_xAddress__reg[9]|Q_net , \cal1_yAddress__reg[0]|Q_net ,
       \cal1_yAddress__reg[10]|Q_net , \cal1_yAddress__reg[1]|Q_net , \cal1_yAddress__reg[2]|Q_net ,
       \cal1_yAddress__reg[3]|Q_net , \cal1_yAddress__reg[4]|Q_net , \cal1_yAddress__reg[5]|Q_net ,
       \cal1_yAddress__reg[6]|Q_net , \cal1_yAddress__reg[7]|Q_net , \cal1_yAddress__reg[8]|Q_net ,
       \cal1_yAddress__reg[9]|Q_net , \coefcal1_divide_inst1_u102_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_10|SUM_net , \coefcal1_divide_inst1_u102_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_12|SUM_net , \coefcal1_divide_inst1_u102_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_14|SUM_net , \coefcal1_divide_inst1_u102_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_1|SUM_net , \coefcal1_divide_inst1_u102_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_3|SUM_net , \coefcal1_divide_inst1_u102_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_5|SUM_net , \coefcal1_divide_inst1_u102_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_7|SUM_net , \coefcal1_divide_inst1_u102_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_9|SUM_net , \coefcal1_divide_inst1_u103_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_10|SUM_net , \coefcal1_divide_inst1_u103_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_12|SUM_net , \coefcal1_divide_inst1_u103_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_14|SUM_net , \coefcal1_divide_inst1_u103_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_1|SUM_net , \coefcal1_divide_inst1_u103_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_3|SUM_net , \coefcal1_divide_inst1_u103_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_5|SUM_net , \coefcal1_divide_inst1_u103_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_7|SUM_net , \coefcal1_divide_inst1_u103_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_9|SUM_net , \coefcal1_divide_inst1_u104_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_10|SUM_net , \coefcal1_divide_inst1_u104_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_12|SUM_net , \coefcal1_divide_inst1_u104_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_14|SUM_net , \coefcal1_divide_inst1_u104_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_1|SUM_net , \coefcal1_divide_inst1_u104_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_3|SUM_net , \coefcal1_divide_inst1_u104_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_5|SUM_net , \coefcal1_divide_inst1_u104_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_7|SUM_net , \coefcal1_divide_inst1_u104_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_9|SUM_net , \coefcal1_divide_inst1_u105_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_10|SUM_net , \coefcal1_divide_inst1_u105_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_12|SUM_net , \coefcal1_divide_inst1_u105_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_14|SUM_net , \coefcal1_divide_inst1_u105_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_1|SUM_net , \coefcal1_divide_inst1_u105_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_3|SUM_net , \coefcal1_divide_inst1_u105_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_5|SUM_net , \coefcal1_divide_inst1_u105_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_7|SUM_net , \coefcal1_divide_inst1_u105_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_9|SUM_net , \coefcal1_divide_inst1_u106_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_10|SUM_net , \coefcal1_divide_inst1_u106_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_12|SUM_net , \coefcal1_divide_inst1_u106_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_14|SUM_net , \coefcal1_divide_inst1_u106_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_1|SUM_net , \coefcal1_divide_inst1_u106_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_3|SUM_net , \coefcal1_divide_inst1_u106_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_5|SUM_net , \coefcal1_divide_inst1_u106_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_7|SUM_net , \coefcal1_divide_inst1_u106_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_9|SUM_net , \coefcal1_divide_inst1_u107_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_10|SUM_net , \coefcal1_divide_inst1_u107_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_12|SUM_net , \coefcal1_divide_inst1_u107_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_14|SUM_net , \coefcal1_divide_inst1_u107_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_1|SUM_net , \coefcal1_divide_inst1_u107_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_3|SUM_net , \coefcal1_divide_inst1_u107_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_5|SUM_net , \coefcal1_divide_inst1_u107_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_7|SUM_net , \coefcal1_divide_inst1_u107_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_9|SUM_net , \coefcal1_divide_inst1_u108_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_10|SUM_net , \coefcal1_divide_inst1_u108_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_12|SUM_net , \coefcal1_divide_inst1_u108_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_14|SUM_net , \coefcal1_divide_inst1_u108_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_1|SUM_net , \coefcal1_divide_inst1_u108_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_3|SUM_net , \coefcal1_divide_inst1_u108_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_5|SUM_net , \coefcal1_divide_inst1_u108_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_7|SUM_net , \coefcal1_divide_inst1_u108_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_9|SUM_net , \coefcal1_divide_inst1_u109_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_10|SUM_net , \coefcal1_divide_inst1_u109_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_12|SUM_net , \coefcal1_divide_inst1_u109_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_14|SUM_net , \coefcal1_divide_inst1_u109_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_1|SUM_net , \coefcal1_divide_inst1_u109_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_3|SUM_net , \coefcal1_divide_inst1_u109_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_5|SUM_net , \coefcal1_divide_inst1_u109_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_7|SUM_net , \coefcal1_divide_inst1_u109_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_9|SUM_net , \coefcal1_divide_inst1_u110_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_10|SUM_net , \coefcal1_divide_inst1_u110_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_12|SUM_net , \coefcal1_divide_inst1_u110_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_14|SUM_net , \coefcal1_divide_inst1_u110_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_1|SUM_net , \coefcal1_divide_inst1_u110_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_3|SUM_net , \coefcal1_divide_inst1_u110_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_5|SUM_net , \coefcal1_divide_inst1_u110_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_7|SUM_net , \coefcal1_divide_inst1_u110_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_9|SUM_net , \coefcal1_divide_inst1_u111_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_10|SUM_net , \coefcal1_divide_inst1_u111_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_12|SUM_net , \coefcal1_divide_inst1_u111_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_14|SUM_net , \coefcal1_divide_inst1_u111_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_1|SUM_net , \coefcal1_divide_inst1_u111_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_3|SUM_net , \coefcal1_divide_inst1_u111_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_5|SUM_net , \coefcal1_divide_inst1_u111_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_7|SUM_net , \coefcal1_divide_inst1_u111_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_9|SUM_net , \coefcal1_divide_inst1_u112_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_10|SUM_net , \coefcal1_divide_inst1_u112_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_12|SUM_net , \coefcal1_divide_inst1_u112_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_14|SUM_net , \coefcal1_divide_inst1_u112_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_1|SUM_net , \coefcal1_divide_inst1_u112_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_3|SUM_net , \coefcal1_divide_inst1_u112_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_5|SUM_net , \coefcal1_divide_inst1_u112_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_7|SUM_net , \coefcal1_divide_inst1_u112_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_9|SUM_net , \coefcal1_divide_inst1_u113_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_10|SUM_net , \coefcal1_divide_inst1_u113_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_12|SUM_net , \coefcal1_divide_inst1_u113_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_14|SUM_net , \coefcal1_divide_inst1_u113_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_1|SUM_net , \coefcal1_divide_inst1_u113_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_3|SUM_net , \coefcal1_divide_inst1_u113_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_5|SUM_net , \coefcal1_divide_inst1_u113_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_7|SUM_net , \coefcal1_divide_inst1_u113_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_9|SUM_net , \coefcal1_divide_inst1_u114_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_10|SUM_net , \coefcal1_divide_inst1_u114_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_12|SUM_net , \coefcal1_divide_inst1_u114_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_14|SUM_net , \coefcal1_divide_inst1_u114_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_1|SUM_net , \coefcal1_divide_inst1_u114_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_3|SUM_net , \coefcal1_divide_inst1_u114_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_5|SUM_net , \coefcal1_divide_inst1_u114_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_7|SUM_net , \coefcal1_divide_inst1_u114_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_9|SUM_net , \coefcal1_divide_inst1_u115_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_10|SUM_net , \coefcal1_divide_inst1_u115_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_12|SUM_net , \coefcal1_divide_inst1_u115_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_14|SUM_net , \coefcal1_divide_inst1_u115_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_1|SUM_net , \coefcal1_divide_inst1_u115_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_3|SUM_net , \coefcal1_divide_inst1_u115_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_5|SUM_net , \coefcal1_divide_inst1_u115_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_7|SUM_net , \coefcal1_divide_inst1_u115_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_9|SUM_net , \coefcal1_divide_inst1_u116_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_10|SUM_net , \coefcal1_divide_inst1_u116_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_12|SUM_net , \coefcal1_divide_inst1_u116_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_14|SUM_net , \coefcal1_divide_inst1_u116_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_1|SUM_net , \coefcal1_divide_inst1_u116_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_3|SUM_net , \coefcal1_divide_inst1_u116_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_5|SUM_net , \coefcal1_divide_inst1_u116_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_7|SUM_net , \coefcal1_divide_inst1_u116_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_9|SUM_net , \coefcal1_divide_inst1_u118_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u120_XORCI_17|SUM_net , \coefcal1_divide_inst1_u122_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u124_XORCI_17|SUM_net , \coefcal1_divide_inst1_u126_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u128_XORCI_17|SUM_net , \coefcal1_divide_inst1_u130_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u132_XORCI_17|SUM_net , \coefcal1_divide_inst1_u134_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u136_XORCI_17|SUM_net , \coefcal1_divide_inst1_u138_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u140_XORCI_17|SUM_net , \coefcal1_divide_inst1_u142_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u144_XORCI_17|SUM_net , \coefcal1_divide_inst1_u146_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u148_XORCI_17|SUM_net , \coefcal1_divide_inst1_u150_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_0|SUM_net , \coefcal1_divide_inst2_u102_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_11|SUM_net , \coefcal1_divide_inst2_u102_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_13|SUM_net , \coefcal1_divide_inst2_u102_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_15|SUM_net , \coefcal1_divide_inst2_u102_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_2|SUM_net , \coefcal1_divide_inst2_u102_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_4|SUM_net , \coefcal1_divide_inst2_u102_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_6|SUM_net , \coefcal1_divide_inst2_u102_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_8|SUM_net , \coefcal1_divide_inst2_u102_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_0|SUM_net , \coefcal1_divide_inst2_u103_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_11|SUM_net , \coefcal1_divide_inst2_u103_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_13|SUM_net , \coefcal1_divide_inst2_u103_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_15|SUM_net , \coefcal1_divide_inst2_u103_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_2|SUM_net , \coefcal1_divide_inst2_u103_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_4|SUM_net , \coefcal1_divide_inst2_u103_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_6|SUM_net , \coefcal1_divide_inst2_u103_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_8|SUM_net , \coefcal1_divide_inst2_u103_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_0|SUM_net , \coefcal1_divide_inst2_u104_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_11|SUM_net , \coefcal1_divide_inst2_u104_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_13|SUM_net , \coefcal1_divide_inst2_u104_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_15|SUM_net , \coefcal1_divide_inst2_u104_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_2|SUM_net , \coefcal1_divide_inst2_u104_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_4|SUM_net , \coefcal1_divide_inst2_u104_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_6|SUM_net , \coefcal1_divide_inst2_u104_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_8|SUM_net , \coefcal1_divide_inst2_u104_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_0|SUM_net , \coefcal1_divide_inst2_u105_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_11|SUM_net , \coefcal1_divide_inst2_u105_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_13|SUM_net , \coefcal1_divide_inst2_u105_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_15|SUM_net , \coefcal1_divide_inst2_u105_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_2|SUM_net , \coefcal1_divide_inst2_u105_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_4|SUM_net , \coefcal1_divide_inst2_u105_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_6|SUM_net , \coefcal1_divide_inst2_u105_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_8|SUM_net , \coefcal1_divide_inst2_u105_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_0|SUM_net , \coefcal1_divide_inst2_u106_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_11|SUM_net , \coefcal1_divide_inst2_u106_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_13|SUM_net , \coefcal1_divide_inst2_u106_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_15|SUM_net , \coefcal1_divide_inst2_u106_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_2|SUM_net , \coefcal1_divide_inst2_u106_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_4|SUM_net , \coefcal1_divide_inst2_u106_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_6|SUM_net , \coefcal1_divide_inst2_u106_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_8|SUM_net , \coefcal1_divide_inst2_u106_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_0|SUM_net , \coefcal1_divide_inst2_u107_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_11|SUM_net , \coefcal1_divide_inst2_u107_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_13|SUM_net , \coefcal1_divide_inst2_u107_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_15|SUM_net , \coefcal1_divide_inst2_u107_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_2|SUM_net , \coefcal1_divide_inst2_u107_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_4|SUM_net , \coefcal1_divide_inst2_u107_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_6|SUM_net , \coefcal1_divide_inst2_u107_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_8|SUM_net , \coefcal1_divide_inst2_u107_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_0|SUM_net , \coefcal1_divide_inst2_u108_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_11|SUM_net , \coefcal1_divide_inst2_u108_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_13|SUM_net , \coefcal1_divide_inst2_u108_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_15|SUM_net , \coefcal1_divide_inst2_u108_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_2|SUM_net , \coefcal1_divide_inst2_u108_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_4|SUM_net , \coefcal1_divide_inst2_u108_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_6|SUM_net , \coefcal1_divide_inst2_u108_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_8|SUM_net , \coefcal1_divide_inst2_u108_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_0|SUM_net , \coefcal1_divide_inst2_u109_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_11|SUM_net , \coefcal1_divide_inst2_u109_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_13|SUM_net , \coefcal1_divide_inst2_u109_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_15|SUM_net , \coefcal1_divide_inst2_u109_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_2|SUM_net , \coefcal1_divide_inst2_u109_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_4|SUM_net , \coefcal1_divide_inst2_u109_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_6|SUM_net , \coefcal1_divide_inst2_u109_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_8|SUM_net , \coefcal1_divide_inst2_u109_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_0|SUM_net , \coefcal1_divide_inst2_u110_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_11|SUM_net , \coefcal1_divide_inst2_u110_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_13|SUM_net , \coefcal1_divide_inst2_u110_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_15|SUM_net , \coefcal1_divide_inst2_u110_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_2|SUM_net , \coefcal1_divide_inst2_u110_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_4|SUM_net , \coefcal1_divide_inst2_u110_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_6|SUM_net , \coefcal1_divide_inst2_u110_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_8|SUM_net , \coefcal1_divide_inst2_u110_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_0|SUM_net , \coefcal1_divide_inst2_u111_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_11|SUM_net , \coefcal1_divide_inst2_u111_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_13|SUM_net , \coefcal1_divide_inst2_u111_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_15|SUM_net , \coefcal1_divide_inst2_u111_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_2|SUM_net , \coefcal1_divide_inst2_u111_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_4|SUM_net , \coefcal1_divide_inst2_u111_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_6|SUM_net , \coefcal1_divide_inst2_u111_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_8|SUM_net , \coefcal1_divide_inst2_u111_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_0|SUM_net , \coefcal1_divide_inst2_u112_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_11|SUM_net , \coefcal1_divide_inst2_u112_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_13|SUM_net , \coefcal1_divide_inst2_u112_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_15|SUM_net , \coefcal1_divide_inst2_u112_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_2|SUM_net , \coefcal1_divide_inst2_u112_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_4|SUM_net , \coefcal1_divide_inst2_u112_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_6|SUM_net , \coefcal1_divide_inst2_u112_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_8|SUM_net , \coefcal1_divide_inst2_u112_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_0|SUM_net , \coefcal1_divide_inst2_u113_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_11|SUM_net , \coefcal1_divide_inst2_u113_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_13|SUM_net , \coefcal1_divide_inst2_u113_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_15|SUM_net , \coefcal1_divide_inst2_u113_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_2|SUM_net , \coefcal1_divide_inst2_u113_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_4|SUM_net , \coefcal1_divide_inst2_u113_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_6|SUM_net , \coefcal1_divide_inst2_u113_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_8|SUM_net , \coefcal1_divide_inst2_u113_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_0|SUM_net , \coefcal1_divide_inst2_u114_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_11|SUM_net , \coefcal1_divide_inst2_u114_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_13|SUM_net , \coefcal1_divide_inst2_u114_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_15|SUM_net , \coefcal1_divide_inst2_u114_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_2|SUM_net , \coefcal1_divide_inst2_u114_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_4|SUM_net , \coefcal1_divide_inst2_u114_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_6|SUM_net , \coefcal1_divide_inst2_u114_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_8|SUM_net , \coefcal1_divide_inst2_u114_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_0|SUM_net , \coefcal1_divide_inst2_u115_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_11|SUM_net , \coefcal1_divide_inst2_u115_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_13|SUM_net , \coefcal1_divide_inst2_u115_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_15|SUM_net , \coefcal1_divide_inst2_u115_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_2|SUM_net , \coefcal1_divide_inst2_u115_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_4|SUM_net , \coefcal1_divide_inst2_u115_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_6|SUM_net , \coefcal1_divide_inst2_u115_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_8|SUM_net , \coefcal1_divide_inst2_u115_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_0|SUM_net , \coefcal1_divide_inst2_u116_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_11|SUM_net , \coefcal1_divide_inst2_u116_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_13|SUM_net , \coefcal1_divide_inst2_u116_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_15|SUM_net , \coefcal1_divide_inst2_u116_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_2|SUM_net , \coefcal1_divide_inst2_u116_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_4|SUM_net , \coefcal1_divide_inst2_u116_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_6|SUM_net , \coefcal1_divide_inst2_u116_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_8|SUM_net , \coefcal1_divide_inst2_u116_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u118_XORCI_17|SUM_net , \coefcal1_divide_inst2_u120_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u122_XORCI_17|SUM_net , \coefcal1_divide_inst2_u124_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u126_XORCI_17|SUM_net , \coefcal1_divide_inst2_u128_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u130_XORCI_17|SUM_net , \coefcal1_divide_inst2_u132_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u134_XORCI_17|SUM_net , \coefcal1_divide_inst2_u136_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u138_XORCI_17|SUM_net , \coefcal1_divide_inst2_u140_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u142_XORCI_17|SUM_net , \coefcal1_divide_inst2_u144_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u146_XORCI_17|SUM_net , \coefcal1_divide_inst2_u148_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u150_XORCI_17|SUM_net , \coefcal1_frameRate__reg[0]|Q_net ,
       \coefcal1_frameRate__reg[1]|Q_net , \coefcal1_frameRate__reg[2]|Q_net ,
       \coefcal1_frameRate__reg[3]|Q_net , \coefcal1_frameRate__reg[4]|Q_net ,
       \coefcal1_frameRate__reg[5]|Q_net , \coefcal1_frameRate__reg[6]|Q_net ,
       \coefcal1_frameRate__reg[7]|Q_net , \coefcal1_frameRate__reg[8]|Q_net ,
       \coefcal1_inEn__reg|Q_net , \coefcal1_u59_XORCI_0|SUM_net , \coefcal1_u59_XORCI_10|SUM_net ,
       \coefcal1_u59_XORCI_1|SUM_net , \coefcal1_u59_XORCI_2|SUM_net , \coefcal1_u59_XORCI_3|SUM_net ,
       \coefcal1_u59_XORCI_4|SUM_net , \coefcal1_u59_XORCI_5|SUM_net , \coefcal1_u59_XORCI_6|SUM_net ,
       \coefcal1_u59_XORCI_7|SUM_net , \coefcal1_u59_XORCI_8|SUM_net , \coefcal1_u59_XORCI_9|SUM_net ,
       \coefcal1_u60_XORCI_0|SUM_net , \coefcal1_u60_XORCI_10|SUM_net , \coefcal1_u60_XORCI_1|SUM_net ,
       \coefcal1_u60_XORCI_2|SUM_net , \coefcal1_u60_XORCI_3|SUM_net , \coefcal1_u60_XORCI_4|SUM_net ,
       \coefcal1_u60_XORCI_5|SUM_net , \coefcal1_u60_XORCI_6|SUM_net , \coefcal1_u60_XORCI_7|SUM_net ,
       \coefcal1_u60_XORCI_8|SUM_net , \coefcal1_u60_XORCI_9|SUM_net , \coefcal1_u61_XORCI_0|SUM_net ,
       \coefcal1_u61_XORCI_1|SUM_net , \coefcal1_u61_XORCI_2|SUM_net , \coefcal1_u61_XORCI_3|SUM_net ,
       \coefcal1_u61_XORCI_4|SUM_net , \coefcal1_u61_XORCI_5|SUM_net , \coefcal1_u61_XORCI_6|SUM_net ,
       \coefcal1_u61_XORCI_7|SUM_net , \coefcal1_u62_XORCI_0|SUM_net , \coefcal1_u62_XORCI_1|SUM_net ,
       \coefcal1_u62_XORCI_2|SUM_net , \coefcal1_u62_XORCI_3|SUM_net , \coefcal1_u62_XORCI_4|SUM_net ,
       \coefcal1_u62_XORCI_5|SUM_net , \coefcal1_u62_XORCI_6|SUM_net , \coefcal1_u62_XORCI_7|SUM_net ,
       \coefcal1_u64_XORCI_0|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , \coefcal1_u64_XORCI_11|SUM_net ,
       \coefcal1_u64_XORCI_12|SUM_net , \coefcal1_u64_XORCI_1|SUM_net , \coefcal1_u64_XORCI_2|SUM_net ,
       \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , \coefcal1_u64_XORCI_5|SUM_net ,
       \coefcal1_u64_XORCI_6|SUM_net , \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_8|SUM_net ,
       \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u7_XORCI_0|SUM_net , \coefcal1_u7_XORCI_10|SUM_net ,
       \coefcal1_u7_XORCI_1|SUM_net , \coefcal1_u7_XORCI_2|SUM_net , \coefcal1_u7_XORCI_3|SUM_net ,
       \coefcal1_u7_XORCI_4|SUM_net , \coefcal1_u7_XORCI_5|SUM_net , \coefcal1_u7_XORCI_6|SUM_net ,
       \coefcal1_u7_XORCI_7|SUM_net , \coefcal1_u7_XORCI_8|SUM_net , \coefcal1_u7_XORCI_9|SUM_net ,
       \coefcal1_u8_XORCI_33|SUM_net , \coefcal1_work__reg|Q_net , \coefcal1_working__reg[0]|Q_net ,
       \coefcal1_working__reg[10]|Q_net , \coefcal1_working__reg[11]|Q_net ,
       \coefcal1_working__reg[12]|Q_net , \coefcal1_working__reg[13]|Q_net ,
       \coefcal1_working__reg[14]|Q_net , \coefcal1_working__reg[15]|Q_net ,
       \coefcal1_working__reg[16]|Q_net , \coefcal1_working__reg[17]|Q_net ,
       \coefcal1_working__reg[18]|Q_net , \coefcal1_working__reg[19]|Q_net ,
       \coefcal1_working__reg[1]|Q_net , \coefcal1_working__reg[20]|Q_net , \coefcal1_working__reg[21]|Q_net ,
       \coefcal1_working__reg[22]|Q_net , \coefcal1_working__reg[23]|Q_net ,
       \coefcal1_working__reg[24]|Q_net , \coefcal1_working__reg[25]|Q_net ,
       \coefcal1_working__reg[26]|Q_net , \coefcal1_working__reg[27]|Q_net ,
       \coefcal1_working__reg[28]|Q_net , \coefcal1_working__reg[29]|Q_net ,
       \coefcal1_working__reg[2]|Q_net , \coefcal1_working__reg[30]|Q_net , \coefcal1_working__reg[31]|Q_net ,
       \coefcal1_working__reg[32]|Q_net , \coefcal1_working__reg[3]|Q_net , \coefcal1_working__reg[4]|Q_net ,
       \coefcal1_working__reg[5]|Q_net , \coefcal1_working__reg[6]|Q_net , \coefcal1_working__reg[7]|Q_net ,
       \coefcal1_working__reg[8]|Q_net , \coefcal1_working__reg[9]|Q_net , \coefcal1_xDividend__reg[0]|Q_net ,
       \coefcal1_xDividend__reg[10]|Q_net , \coefcal1_xDividend__reg[11]|Q_net ,
       \coefcal1_xDividend__reg[12]|Q_net , \coefcal1_xDividend__reg[13]|Q_net ,
       \coefcal1_xDividend__reg[14]|Q_net , \coefcal1_xDividend__reg[15]|Q_net ,
       \coefcal1_xDividend__reg[16]|Q_net , \coefcal1_xDividend__reg[1]|Q_net ,
       \coefcal1_xDividend__reg[2]|Q_net , \coefcal1_xDividend__reg[3]|Q_net ,
       \coefcal1_xDividend__reg[4]|Q_net , \coefcal1_xDividend__reg[5]|Q_net ,
       \coefcal1_xDividend__reg[6]|Q_net , \coefcal1_xDividend__reg[7]|Q_net ,
       \coefcal1_xDividend__reg[8]|Q_net , \coefcal1_xDividend__reg[9]|Q_net ,
       \coefcal1_xDivisor__reg[0]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net ,
       \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net ,
       \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net ,
       \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[16]|Q_net ,
       \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net ,
       \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net ,
       \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net ,
       \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net ,
       \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_yDividend__reg[0]|Q_net ,
       \coefcal1_yDividend__reg[10]|Q_net , \coefcal1_yDividend__reg[11]|Q_net ,
       \coefcal1_yDividend__reg[12]|Q_net , \coefcal1_yDividend__reg[13]|Q_net ,
       \coefcal1_yDividend__reg[14]|Q_net , \coefcal1_yDividend__reg[15]|Q_net ,
       \coefcal1_yDividend__reg[16]|Q_net , \coefcal1_yDividend__reg[1]|Q_net ,
       \coefcal1_yDividend__reg[2]|Q_net , \coefcal1_yDividend__reg[3]|Q_net ,
       \coefcal1_yDividend__reg[4]|Q_net , \coefcal1_yDividend__reg[5]|Q_net ,
       \coefcal1_yDividend__reg[6]|Q_net , \coefcal1_yDividend__reg[7]|Q_net ,
       \coefcal1_yDividend__reg[8]|Q_net , \coefcal1_yDividend__reg[9]|Q_net ,
       \coefcal1_yDivisor__reg[0]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net ,
       \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net ,
       \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net ,
       \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[16]|Q_net ,
       \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net ,
       \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net ,
       \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net ,
       \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net ,
       \coefcal1_yDivisor__reg[9]|Q_net , \fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_0_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_1_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_1_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_3_ab_reg__reg[0]|Q_net , \inputctrl1_dataOut__reg[0]|Q_net ,
       \inputctrl1_dataOut__reg[10]|Q_net , \inputctrl1_dataOut__reg[11]|Q_net ,
       \inputctrl1_dataOut__reg[12]|Q_net , \inputctrl1_dataOut__reg[13]|Q_net ,
       \inputctrl1_dataOut__reg[14]|Q_net , \inputctrl1_dataOut__reg[15]|Q_net ,
       \inputctrl1_dataOut__reg[1]|Q_net , \inputctrl1_dataOut__reg[2]|Q_net ,
       \inputctrl1_dataOut__reg[3]|Q_net , \inputctrl1_dataOut__reg[4]|Q_net ,
       \inputctrl1_dataOut__reg[5]|Q_net , \inputctrl1_dataOut__reg[6]|Q_net ,
       \inputctrl1_dataOut__reg[7]|Q_net , \inputctrl1_dataOut__reg[8]|Q_net ,
       \inputctrl1_dataOut__reg[9]|Q_net , \inputctrl1_jmp__reg|Q_net , \inputctrl1_ramWrtAddr__reg[0]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[10]|Q_net , \inputctrl1_ramWrtAddr__reg[1]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[2]|Q_net , \inputctrl1_ramWrtAddr__reg[3]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[4]|Q_net , \inputctrl1_ramWrtAddr__reg[5]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[6]|Q_net , \inputctrl1_ramWrtAddr__reg[7]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[8]|Q_net , \inputctrl1_ramWrtAddr__reg[9]|Q_net ,
       \inputctrl1_ramWrtEn__reg|Q_net , \inputctrl1_u108_XORCI_0|SUM_net , \inputctrl1_u108_XORCI_10|SUM_net ,
       \inputctrl1_u108_XORCI_11|SUM_net , \inputctrl1_u108_XORCI_12|SUM_net ,
       \inputctrl1_u108_XORCI_13|SUM_net , \inputctrl1_u108_XORCI_14|SUM_net ,
       \inputctrl1_u108_XORCI_15|SUM_net , \inputctrl1_u108_XORCI_16|SUM_net ,
       \inputctrl1_u108_XORCI_1|SUM_net , \inputctrl1_u108_XORCI_2|SUM_net ,
       \inputctrl1_u108_XORCI_3|SUM_net , \inputctrl1_u108_XORCI_4|SUM_net ,
       \inputctrl1_u108_XORCI_5|SUM_net , \inputctrl1_u108_XORCI_6|SUM_net ,
       \inputctrl1_u108_XORCI_7|SUM_net , \inputctrl1_u108_XORCI_8|SUM_net ,
       \inputctrl1_u108_XORCI_9|SUM_net , \inputctrl1_u109_XORCI_0|SUM_net ,
       \inputctrl1_u109_XORCI_10|SUM_net , \inputctrl1_u109_XORCI_11|SUM_net ,
       \inputctrl1_u109_XORCI_12|SUM_net , \inputctrl1_u109_XORCI_13|SUM_net ,
       \inputctrl1_u109_XORCI_14|SUM_net , \inputctrl1_u109_XORCI_15|SUM_net ,
       \inputctrl1_u109_XORCI_16|SUM_net , \inputctrl1_u109_XORCI_1|SUM_net ,
       \inputctrl1_u109_XORCI_2|SUM_net , \inputctrl1_u109_XORCI_3|SUM_net ,
       \inputctrl1_u109_XORCI_4|SUM_net , \inputctrl1_u109_XORCI_5|SUM_net ,
       \inputctrl1_u109_XORCI_6|SUM_net , \inputctrl1_u109_XORCI_7|SUM_net ,
       \inputctrl1_u109_XORCI_8|SUM_net , \inputctrl1_u109_XORCI_9|SUM_net ,
       \inputctrl1_u110_XORCI_0|SUM_net , \inputctrl1_u110_XORCI_10|SUM_net ,
       \inputctrl1_u110_XORCI_1|SUM_net , \inputctrl1_u110_XORCI_2|SUM_net ,
       \inputctrl1_u110_XORCI_3|SUM_net , \inputctrl1_u110_XORCI_4|SUM_net ,
       \inputctrl1_u110_XORCI_5|SUM_net , \inputctrl1_u110_XORCI_6|SUM_net ,
       \inputctrl1_u110_XORCI_7|SUM_net , \inputctrl1_u110_XORCI_8|SUM_net ,
       \inputctrl1_u110_XORCI_9|SUM_net , \inputctrl1_u111_XORCI_0|SUM_net ,
       \inputctrl1_u111_XORCI_10|SUM_net , \inputctrl1_u111_XORCI_1|SUM_net ,
       \inputctrl1_u111_XORCI_2|SUM_net , \inputctrl1_u111_XORCI_3|SUM_net ,
       \inputctrl1_u111_XORCI_4|SUM_net , \inputctrl1_u111_XORCI_5|SUM_net ,
       \inputctrl1_u111_XORCI_6|SUM_net , \inputctrl1_u111_XORCI_7|SUM_net ,
       \inputctrl1_u111_XORCI_8|SUM_net , \inputctrl1_u111_XORCI_9|SUM_net ,
       \inputctrl1_u112_XORCI_0|SUM_net , \inputctrl1_u112_XORCI_10|SUM_net ,
       \inputctrl1_u112_XORCI_1|SUM_net , \inputctrl1_u112_XORCI_2|SUM_net ,
       \inputctrl1_u112_XORCI_3|SUM_net , \inputctrl1_u112_XORCI_4|SUM_net ,
       \inputctrl1_u112_XORCI_5|SUM_net , \inputctrl1_u112_XORCI_6|SUM_net ,
       \inputctrl1_u112_XORCI_7|SUM_net , \inputctrl1_u112_XORCI_8|SUM_net ,
       \inputctrl1_u112_XORCI_9|SUM_net , \inputctrl1_u37_XORCI_11|SUM_net ,
       \inputctrl1_u39_XORCI_11|SUM_net , \inputctrl1_u41_XORCI_11|SUM_net ,
       \inputctrl1_u43_XORCI_11|SUM_net , \inputctrl1_xAddress__reg[0]|Q_net ,
       \inputctrl1_xAddress__reg[10]|Q_net , \inputctrl1_xAddress__reg[1]|Q_net ,
       \inputctrl1_xAddress__reg[2]|Q_net , \inputctrl1_xAddress__reg[3]|Q_net ,
       \inputctrl1_xAddress__reg[4]|Q_net , \inputctrl1_xAddress__reg[5]|Q_net ,
       \inputctrl1_xAddress__reg[6]|Q_net , \inputctrl1_xAddress__reg[7]|Q_net ,
       \inputctrl1_xAddress__reg[8]|Q_net , \inputctrl1_xAddress__reg[9]|Q_net ,
       \inputctrl1_xCal__reg[0]|Q_net , \inputctrl1_xCal__reg[10]|Q_net , \inputctrl1_xCal__reg[11]|Q_net ,
       \inputctrl1_xCal__reg[12]|Q_net , \inputctrl1_xCal__reg[13]|Q_net , \inputctrl1_xCal__reg[14]|Q_net ,
       \inputctrl1_xCal__reg[15]|Q_net , \inputctrl1_xCal__reg[16]|Q_net , \inputctrl1_xCal__reg[1]|Q_net ,
       \inputctrl1_xCal__reg[2]|Q_net , \inputctrl1_xCal__reg[3]|Q_net , \inputctrl1_xCal__reg[4]|Q_net ,
       \inputctrl1_xCal__reg[5]|Q_net , \inputctrl1_xCal__reg[6]|Q_net , \inputctrl1_xCal__reg[7]|Q_net ,
       \inputctrl1_xCal__reg[8]|Q_net , \inputctrl1_xCal__reg[9]|Q_net , \inputctrl1_xPreEn__reg|Q_net ,
       \inputctrl1_yAddress__reg[0]|Q_net , \inputctrl1_yAddress__reg[10]|Q_net ,
       \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net ,
       \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net ,
       \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net ,
       \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net ,
       \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yCal__reg[0]|Q_net ,
       \inputctrl1_yCal__reg[10]|Q_net , \inputctrl1_yCal__reg[11]|Q_net , \inputctrl1_yCal__reg[12]|Q_net ,
       \inputctrl1_yCal__reg[13]|Q_net , \inputctrl1_yCal__reg[14]|Q_net , \inputctrl1_yCal__reg[15]|Q_net ,
       \inputctrl1_yCal__reg[16]|Q_net , \inputctrl1_yCal__reg[1]|Q_net , \inputctrl1_yCal__reg[2]|Q_net ,
       \inputctrl1_yCal__reg[3]|Q_net , \inputctrl1_yCal__reg[4]|Q_net , \inputctrl1_yCal__reg[5]|Q_net ,
       \inputctrl1_yCal__reg[6]|Q_net , \inputctrl1_yCal__reg[7]|Q_net , \inputctrl1_yCal__reg[8]|Q_net ,
       \inputctrl1_yCal__reg[9]|Q_net , \inputctrl1_yPreEn__reg|Q_net , \u2_XORCI_0|SUM_net ,
       \u2_XORCI_10|SUM_net , \u2_XORCI_11|SUM_net , \u2_XORCI_1|SUM_net , \u2_XORCI_2|SUM_net ,
       \u2_XORCI_3|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_5|SUM_net , \u2_XORCI_6|SUM_net ,
       \u2_XORCI_7|SUM_net , \u2_XORCI_8|SUM_net , \u2_XORCI_9|SUM_net , \u3_XORCI_0|SUM_net ,
       \u3_XORCI_10|SUM_net , \u3_XORCI_1|SUM_net , \u3_XORCI_2|SUM_net , \u3_XORCI_3|SUM_net ,
       \u3_XORCI_4|SUM_net , \u3_XORCI_5|SUM_net , \u3_XORCI_6|SUM_net , \u3_XORCI_7|SUM_net ,
       \u3_XORCI_8|SUM_net , \u3_XORCI_9|SUM_net ;

    assign HS = HS_1863_net;
    assign a_acc_en_cal1_u135_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u136_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u137_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u138_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u139_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u140_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u141_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u142_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u143_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u144_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u145_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_cal1_u146_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_coefcal1_u63_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign a_acc_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign \a_dinx[0]_cal1_u134_mac  = \cal1_uPreF__reg[0]|Q_net ;
    assign \a_dinx[0]_cal1_u135_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_dinx[0]_cal1_u138_mac  = \a_mac_out[6]_cal1_u134_mac ;
    assign \a_dinx[0]_cal1_u139_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_dinx[0]_cal1_u140_mac  = \a_dinx[0]_cal1_u136_mac ;
    assign \a_dinx[0]_cal1_u141_mac  = \a_dinx[0]_cal1_u137_mac ;
    assign \a_dinx[0]_cal1_u142_mac  = \a_mac_out[6]_cal1_u134_mac ;
    assign \a_dinx[0]_cal1_u143_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_dinx[0]_cal1_u144_mac  = \a_dinx[0]_cal1_u136_mac ;
    assign \a_dinx[0]_cal1_u145_mac  = \a_dinx[0]_cal1_u137_mac ;
    assign \a_dinx[0]_cal1_u146_mac  = \a_mac_out[6]_cal1_u134_mac ;
    assign \a_dinx[0]_coefcal1_u63_mac  = outYRes[0];
    assign \a_dinx[0]_coefcal1_u64_mac  = \a_mac_out[0]_coefcal1_u63_mac ;
    assign \a_dinx[0]_coefcal1_u64_mac_0_  = \a_mac_out[18]_coefcal1_u63_mac ;
    assign \a_dinx[10]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_coefcal1_u63_mac  = outYRes[10];
    assign \a_dinx[10]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[10]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_coefcal1_u63_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[11]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_coefcal1_u63_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[12]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_coefcal1_u63_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[13]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[1]_cal1_u134_mac  = \cal1_uPreF__reg[1]|Q_net ;
    assign \a_dinx[1]_cal1_u135_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_dinx[1]_cal1_u138_mac  = \a_mac_out[7]_cal1_u134_mac ;
    assign \a_dinx[1]_cal1_u139_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_dinx[1]_cal1_u140_mac  = \a_dinx[1]_cal1_u136_mac ;
    assign \a_dinx[1]_cal1_u141_mac  = \a_dinx[1]_cal1_u137_mac ;
    assign \a_dinx[1]_cal1_u142_mac  = \a_mac_out[7]_cal1_u134_mac ;
    assign \a_dinx[1]_cal1_u143_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_dinx[1]_cal1_u144_mac  = \a_dinx[1]_cal1_u136_mac ;
    assign \a_dinx[1]_cal1_u145_mac  = \a_dinx[1]_cal1_u137_mac ;
    assign \a_dinx[1]_cal1_u146_mac  = \a_mac_out[7]_cal1_u134_mac ;
    assign \a_dinx[1]_coefcal1_u63_mac  = outYRes[1];
    assign \a_dinx[1]_coefcal1_u64_mac  = \a_mac_out[1]_coefcal1_u63_mac ;
    assign \a_dinx[1]_coefcal1_u64_mac_0_  = \a_mac_out[19]_coefcal1_u63_mac ;
    assign \a_dinx[2]_cal1_u134_mac  = \cal1_uPreF__reg[2]|Q_net ;
    assign \a_dinx[2]_cal1_u135_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_dinx[2]_cal1_u138_mac  = \a_mac_out[8]_cal1_u134_mac ;
    assign \a_dinx[2]_cal1_u139_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_dinx[2]_cal1_u140_mac  = \a_dinx[2]_cal1_u136_mac ;
    assign \a_dinx[2]_cal1_u141_mac  = \a_dinx[2]_cal1_u137_mac ;
    assign \a_dinx[2]_cal1_u142_mac  = \a_mac_out[8]_cal1_u134_mac ;
    assign \a_dinx[2]_cal1_u143_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_dinx[2]_cal1_u144_mac  = \a_dinx[2]_cal1_u136_mac ;
    assign \a_dinx[2]_cal1_u145_mac  = \a_dinx[2]_cal1_u137_mac ;
    assign \a_dinx[2]_cal1_u146_mac  = \a_mac_out[8]_cal1_u134_mac ;
    assign \a_dinx[2]_coefcal1_u63_mac  = outYRes[2];
    assign \a_dinx[2]_coefcal1_u64_mac  = \a_mac_out[2]_coefcal1_u63_mac ;
    assign \a_dinx[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[3]_cal1_u134_mac  = \cal1_uPreF__reg[3]|Q_net ;
    assign \a_dinx[3]_cal1_u135_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_dinx[3]_cal1_u138_mac  = \a_mac_out[9]_cal1_u134_mac ;
    assign \a_dinx[3]_cal1_u139_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_dinx[3]_cal1_u140_mac  = \a_dinx[3]_cal1_u136_mac ;
    assign \a_dinx[3]_cal1_u141_mac  = \a_dinx[3]_cal1_u137_mac ;
    assign \a_dinx[3]_cal1_u142_mac  = \a_mac_out[9]_cal1_u134_mac ;
    assign \a_dinx[3]_cal1_u143_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_dinx[3]_cal1_u144_mac  = \a_dinx[3]_cal1_u136_mac ;
    assign \a_dinx[3]_cal1_u145_mac  = \a_dinx[3]_cal1_u137_mac ;
    assign \a_dinx[3]_cal1_u146_mac  = \a_mac_out[9]_cal1_u134_mac ;
    assign \a_dinx[3]_coefcal1_u63_mac  = outYRes[3];
    assign \a_dinx[3]_coefcal1_u64_mac  = \a_mac_out[3]_coefcal1_u63_mac ;
    assign \a_dinx[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[4]_cal1_u134_mac  = \cal1_uPreF__reg[4]|Q_net ;
    assign \a_dinx[4]_cal1_u135_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_dinx[4]_cal1_u138_mac  = \a_mac_out[10]_cal1_u134_mac ;
    assign \a_dinx[4]_cal1_u139_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_dinx[4]_cal1_u140_mac  = \a_dinx[4]_cal1_u136_mac ;
    assign \a_dinx[4]_cal1_u141_mac  = \a_dinx[4]_cal1_u137_mac ;
    assign \a_dinx[4]_cal1_u142_mac  = \a_mac_out[10]_cal1_u134_mac ;
    assign \a_dinx[4]_cal1_u143_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_dinx[4]_cal1_u144_mac  = \a_dinx[4]_cal1_u136_mac ;
    assign \a_dinx[4]_cal1_u145_mac  = \a_dinx[4]_cal1_u137_mac ;
    assign \a_dinx[4]_cal1_u146_mac  = \a_mac_out[10]_cal1_u134_mac ;
    assign \a_dinx[4]_coefcal1_u63_mac  = outYRes[4];
    assign \a_dinx[4]_coefcal1_u64_mac  = \a_mac_out[4]_coefcal1_u63_mac ;
    assign \a_dinx[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[5]_cal1_u134_mac  = \cal1_uPreF__reg[5]|Q_net ;
    assign \a_dinx[5]_cal1_u135_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_dinx[5]_cal1_u138_mac  = \a_mac_out[11]_cal1_u134_mac ;
    assign \a_dinx[5]_cal1_u139_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_dinx[5]_cal1_u140_mac  = \a_dinx[5]_cal1_u136_mac ;
    assign \a_dinx[5]_cal1_u141_mac  = \a_dinx[5]_cal1_u137_mac ;
    assign \a_dinx[5]_cal1_u142_mac  = \a_mac_out[11]_cal1_u134_mac ;
    assign \a_dinx[5]_cal1_u143_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_dinx[5]_cal1_u144_mac  = \a_dinx[5]_cal1_u136_mac ;
    assign \a_dinx[5]_cal1_u145_mac  = \a_dinx[5]_cal1_u137_mac ;
    assign \a_dinx[5]_cal1_u146_mac  = \a_mac_out[11]_cal1_u134_mac ;
    assign \a_dinx[5]_coefcal1_u63_mac  = outYRes[5];
    assign \a_dinx[5]_coefcal1_u64_mac  = \a_mac_out[5]_coefcal1_u63_mac ;
    assign \a_dinx[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u135_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_dinx[6]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u139_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_dinx[6]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u143_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_dinx[6]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_coefcal1_u63_mac  = outYRes[6];
    assign \a_dinx[6]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_coefcal1_u63_mac  = outYRes[7];
    assign \a_dinx[7]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_coefcal1_u63_mac  = outYRes[8];
    assign \a_dinx[8]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_coefcal1_u63_mac  = outYRes[9];
    assign \a_dinx[9]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_dinx[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u135_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u136_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u137_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u138_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u139_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u140_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u141_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u142_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u143_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u144_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u145_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_cal1_u146_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinxy_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign \a_diny[0]_cal1_u134_mac  = \cal1_v__reg[0]|Q_net ;
    assign \a_diny[0]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[0]|Q_net ;
    assign \a_diny[0]_coefcal1_u64_mac  = outXRes[0];
    assign \a_diny[0]_coefcal1_u64_mac_0_  = outXRes[0];
    assign \a_diny[1]_cal1_u134_mac  = \cal1_v__reg[1]|Q_net ;
    assign \a_diny[1]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[1]|Q_net ;
    assign \a_diny[1]_coefcal1_u64_mac  = outXRes[1];
    assign \a_diny[1]_coefcal1_u64_mac_0_  = outXRes[1];
    assign \a_diny[2]_cal1_u134_mac  = \cal1_v__reg[2]|Q_net ;
    assign \a_diny[2]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[2]|Q_net ;
    assign \a_diny[2]_coefcal1_u64_mac  = outXRes[2];
    assign \a_diny[2]_coefcal1_u64_mac_0_  = outXRes[2];
    assign \a_diny[3]_cal1_u134_mac  = \cal1_v__reg[3]|Q_net ;
    assign \a_diny[3]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[3]|Q_net ;
    assign \a_diny[3]_coefcal1_u64_mac  = outXRes[3];
    assign \a_diny[3]_coefcal1_u64_mac_0_  = outXRes[3];
    assign \a_diny[4]_cal1_u134_mac  = \cal1_v__reg[4]|Q_net ;
    assign \a_diny[4]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[4]|Q_net ;
    assign \a_diny[4]_coefcal1_u64_mac  = outXRes[4];
    assign \a_diny[4]_coefcal1_u64_mac_0_  = outXRes[4];
    assign \a_diny[5]_cal1_u134_mac  = \cal1_v__reg[5]|Q_net ;
    assign \a_diny[5]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[5]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[5]|Q_net ;
    assign \a_diny[5]_coefcal1_u64_mac  = outXRes[5];
    assign \a_diny[5]_coefcal1_u64_mac_0_  = outXRes[5];
    assign \a_diny[6]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[6]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[6]|Q_net ;
    assign \a_diny[6]_coefcal1_u64_mac  = outXRes[6];
    assign \a_diny[6]_coefcal1_u64_mac_0_  = outXRes[6];
    assign \a_diny[7]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[7]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[7]|Q_net ;
    assign \a_diny[7]_coefcal1_u64_mac  = outXRes[7];
    assign \a_diny[7]_coefcal1_u64_mac_0_  = outXRes[7];
    assign \a_diny[8]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[8]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[8]|Q_net ;
    assign \a_diny[8]_coefcal1_u64_mac  = outXRes[8];
    assign \a_diny[8]_coefcal1_u64_mac_0_  = outXRes[8];
    assign \a_diny[9]_cal1_u134_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u135_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u136_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u137_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u138_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u139_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u140_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u141_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u142_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u143_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u144_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u145_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_cal1_u146_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_coefcal1_u63_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \a_diny[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign a_dinz_cen_cal1_u134_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u135_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u136_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u137_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u138_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u139_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u140_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u141_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u142_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u143_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u144_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u145_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_cal1_u146_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign a_dinz_en_cal1_u134_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u135_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u136_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u137_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u138_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u139_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u140_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u141_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u142_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u143_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u144_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u145_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_cal1_u146_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_coefcal1_u63_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign a_dinz_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign a_in_sr_cal1_u134_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u135_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u136_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u137_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u138_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u139_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u140_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u141_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u142_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u143_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u144_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u145_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_cal1_u146_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_coefcal1_u63_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_in_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u134_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u135_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u136_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u137_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u138_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u139_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u140_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u141_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u142_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u143_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u144_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u145_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_cal1_u146_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_mac_out_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u134_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u135_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u136_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u137_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u138_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u139_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u140_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u141_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u142_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u143_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u144_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u145_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_cal1_u146_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_coefcal1_u63_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign a_out_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign a_sload_cal1_u134_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u135_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u136_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u137_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u138_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u139_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u140_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u141_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u142_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u143_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u144_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u145_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_cal1_u146_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_coefcal1_u63_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign a_sload_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign b_acc_en_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign b_acc_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign \b_dinx[0]_coefcal1_u64_mac  = \a_mac_out[6]_coefcal1_u63_mac ;
    assign \b_dinx[0]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[10]_coefcal1_u64_mac  = \a_mac_out[16]_coefcal1_u63_mac ;
    assign \b_dinx[10]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[11]_coefcal1_u64_mac  = \a_mac_out[17]_coefcal1_u63_mac ;
    assign \b_dinx[11]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[12]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[12]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[13]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[13]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[1]_coefcal1_u64_mac  = \a_mac_out[7]_coefcal1_u63_mac ;
    assign \b_dinx[1]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[2]_coefcal1_u64_mac  = \a_mac_out[8]_coefcal1_u63_mac ;
    assign \b_dinx[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[3]_coefcal1_u64_mac  = \a_mac_out[9]_coefcal1_u63_mac ;
    assign \b_dinx[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[4]_coefcal1_u64_mac  = \a_mac_out[10]_coefcal1_u63_mac ;
    assign \b_dinx[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[5]_coefcal1_u64_mac  = \a_mac_out[11]_coefcal1_u63_mac ;
    assign \b_dinx[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[6]_coefcal1_u64_mac  = \a_mac_out[12]_coefcal1_u63_mac ;
    assign \b_dinx[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[7]_coefcal1_u64_mac  = \a_mac_out[13]_coefcal1_u63_mac ;
    assign \b_dinx[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[8]_coefcal1_u64_mac  = \a_mac_out[14]_coefcal1_u63_mac ;
    assign \b_dinx[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_dinx[9]_coefcal1_u64_mac  = \a_mac_out[15]_coefcal1_u63_mac ;
    assign \b_dinx[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign b_dinxy_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign b_dinxy_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign \b_diny[0]_coefcal1_u64_mac  = outXRes[9];
    assign \b_diny[0]_coefcal1_u64_mac_0_  = outXRes[9];
    assign \b_diny[1]_coefcal1_u64_mac  = outXRes[10];
    assign \b_diny[1]_coefcal1_u64_mac_0_  = outXRes[10];
    assign \b_diny[2]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[3]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[4]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[5]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[6]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[7]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[8]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign \b_diny[9]_coefcal1_u64_mac  = a_acc_en_cal1_u134_mac;
    assign \b_diny[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u134_mac;
    assign b_dinz_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign b_dinz_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign b_dinz_en_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign b_dinz_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign b_in_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign b_in_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign b_mac_out_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign b_mac_out_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign b_out_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u134_mac;
    assign b_out_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u134_mac;
    assign b_sload_coefcal1_u64_mac = a_acc_en_cal1_u134_mac;
    assign b_sload_coefcal1_u64_mac_0_ = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign c1r1_clka_fifo1_ram_inst_0_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_1_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r1_clkb_fifo1_ram_inst_0_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_0_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3_u_emb18k_1 = clkb;
    assign \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstna_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_clka_fifo1_ram_inst_0_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_0_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r2_clkb_fifo1_ram_inst_0_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_0_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3_u_emb18k_1 = clkb;
    assign \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstna_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_clka_fifo1_ram_inst_0_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_0_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r3_clkb_fifo1_ram_inst_0_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_0_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3_u_emb18k_1 = clkb;
    assign \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstna_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_clka_fifo1_ram_inst_0_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_0_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1_u_emb18k_0;
    assign c1r4_clkb_fifo1_ram_inst_0_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_0_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3_u_emb18k_1 = clkb;
    assign \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_0_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_1_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_2_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_0  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_3_u_emb18k_1  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstna_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign cea_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_0_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_0_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_1_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_1_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_2_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_2_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_3_u_emb18k_0 = a_dinxy_cen_cal1_u134_mac;
    assign ceb_fifo1_ram_inst_3_u_emb18k_1 = a_dinxy_cen_cal1_u134_mac;
    assign \haa[0]_fifo1_ram_inst_0_u_emb18k_1  = \haa[0]_fifo1_ram_inst_0_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_1_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_2_u_emb18k_1  = \haa[0]_fifo1_ram_inst_2_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1_u_emb18k_0 ;
    assign \haa[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \haa[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \hab[0]_fifo1_ram_inst_0_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_0_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[1]_fifo1_ram_inst_0_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_0_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_1_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_1_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_2_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_2_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_3_u_emb18k_0  = a_acc_en_cal1_u134_mac;
    assign \hab[1]_fifo1_ram_inst_3_u_emb18k_1  = a_acc_en_cal1_u134_mac;
    assign u3662_O_4_ = u3662_O;
    assign u6776_O_1_ = u6776_O;
    assign u6776_O_2_ = u6776_O;
    assign wea_fifo1_ram_inst_0_u_emb18k_1 = wea_fifo1_ram_inst_0_u_emb18k_0;
    assign wea_fifo1_ram_inst_1_u_emb18k_1 = wea_fifo1_ram_inst_1_u_emb18k_0;
    assign wea_fifo1_ram_inst_2_u_emb18k_0 = wea_fifo1_ram_inst_1_u_emb18k_0;
    assign wea_fifo1_ram_inst_2_u_emb18k_1 = wea_fifo1_ram_inst_1_u_emb18k_0;
    assign wea_fifo1_ram_inst_3_u_emb18k_0 = wea_fifo1_ram_inst_1_u_emb18k_0;
    assign wea_fifo1_ram_inst_3_u_emb18k_1 = wea_fifo1_ram_inst_1_u_emb18k_0;
    assign web_fifo1_ram_inst_0_u_emb18k_0 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_0_u_emb18k_1 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_1_u_emb18k_0 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_1_u_emb18k_1 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_2_u_emb18k_0 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_2_u_emb18k_1 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_3_u_emb18k_0 = a_acc_en_cal1_u134_mac;
    assign web_fifo1_ram_inst_3_u_emb18k_1 = a_acc_en_cal1_u134_mac;

    CS_LUT4_PRIM ii0730 ( .DX(VS), .F0(\cal1_VSNormal__reg|Q_net ), .F1(\cal1_enforceJmp__reg|Q_net ), .F2(dummy_abc_1_), .F3(dummy_abc_2_) );
      defparam ii0730.CONFIG_DATA = 16'hEEEE;
      defparam ii0730.PLACE_LOCATION = "NONE";
      defparam ii0730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0731 ( .DX(a_acc_en_cal1_u134_mac), .F0(dummy_abc_3_), .F1(dummy_abc_4_), .F2(dummy_abc_5_), .F3(dummy_abc_6_) );
      defparam ii0731.CONFIG_DATA = 16'h0000;
      defparam ii0731.PLACE_LOCATION = "NONE";
      defparam ii0731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0732 ( .DX(nn0732), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[0]|Q_net ), .F2(\cal1_v__reg[0]|Q_net ), .F3(dummy_abc_7_) );
      defparam ii0732.CONFIG_DATA = 16'h9696;
      defparam ii0732.PLACE_LOCATION = "NONE";
      defparam ii0732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0733 ( .DX(a_dinxy_cen_cal1_u134_mac), .F0(dummy_abc_8_), .F1(dummy_abc_9_), .F2(dummy_abc_10_), .F3(dummy_abc_11_) );
      defparam ii0733.CONFIG_DATA = 16'hFFFF;
      defparam ii0733.PLACE_LOCATION = "NONE";
      defparam ii0733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0734 ( .DX(nn0734), .F0(\cal1_uPreF__reg[0]|Q_net ), .F1(dummy_abc_12_), .F2(dummy_abc_13_), .F3(dummy_abc_14_) );
      defparam ii0734.CONFIG_DATA = 16'h5555;
      defparam ii0734.PLACE_LOCATION = "NONE";
      defparam ii0734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0735 ( .DX(nn0735), .F0(\cal1_uPreF__reg[1]|Q_net ), .F1(dummy_abc_15_), .F2(dummy_abc_16_), .F3(dummy_abc_17_) );
      defparam ii0735.CONFIG_DATA = 16'h5555;
      defparam ii0735.PLACE_LOCATION = "NONE";
      defparam ii0735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0736 ( .DX(nn0736), .F0(\cal1_uPreF__reg[2]|Q_net ), .F1(dummy_abc_18_), .F2(dummy_abc_19_), .F3(dummy_abc_20_) );
      defparam ii0736.CONFIG_DATA = 16'h5555;
      defparam ii0736.PLACE_LOCATION = "NONE";
      defparam ii0736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0737 ( .DX(nn0737), .F0(\cal1_uPreF__reg[3]|Q_net ), .F1(dummy_abc_21_), .F2(dummy_abc_22_), .F3(dummy_abc_23_) );
      defparam ii0737.CONFIG_DATA = 16'h5555;
      defparam ii0737.PLACE_LOCATION = "NONE";
      defparam ii0737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0738 ( .DX(nn0738), .F0(\cal1_uPreF__reg[4]|Q_net ), .F1(dummy_abc_24_), .F2(dummy_abc_25_), .F3(dummy_abc_26_) );
      defparam ii0738.CONFIG_DATA = 16'h5555;
      defparam ii0738.PLACE_LOCATION = "NONE";
      defparam ii0738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0739 ( .DX(nn0739), .F0(\cal1_uPreF__reg[5]|Q_net ), .F1(dummy_abc_27_), .F2(dummy_abc_28_), .F3(dummy_abc_29_) );
      defparam ii0739.CONFIG_DATA = 16'h5555;
      defparam ii0739.PLACE_LOCATION = "NONE";
      defparam ii0739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0740 ( .DX(nn0740), .F0(dummy_abc_30_), .F1(dummy_abc_31_), .F2(dummy_abc_32_), .F3(dummy_abc_33_) );
      defparam ii0740.CONFIG_DATA = 16'h0000;
      defparam ii0740.PLACE_LOCATION = "NONE";
      defparam ii0740.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7_4_ ( 
        .CA( {a_dinxy_cen_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_884_ ), 
        .DX( {nn0740, nn0739, nn0738, nn0737, nn0736, nn0735, nn0734} ), 
        .SUM( {\cal1_u54_XORCI_6|SUM_net , \cal1_u54_XORCI_5|SUM_net , 
              \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_3|SUM_net , \cal1_u54_XORCI_2|SUM_net , 
              \cal1_u54_XORCI_1|SUM_net , \cal1_u54_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0750 ( .DX(nn0750), .F0(\cal1_uPreF__reg[0]|Q_net ), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_abc_34_), .F3(dummy_abc_35_) );
      defparam ii0750.CONFIG_DATA = 16'h9999;
      defparam ii0750.PLACE_LOCATION = "NONE";
      defparam ii0750.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0751 ( .DX(nn0751), .F0(\cal1_v__reg[1]|Q_net ), .F1(\cal1_u54_XORCI_1|SUM_net ), .F2(dummy_abc_36_), .F3(dummy_abc_37_) );
      defparam ii0751.CONFIG_DATA = 16'h9999;
      defparam ii0751.PLACE_LOCATION = "NONE";
      defparam ii0751.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0752 ( .DX(nn0752), .F0(\cal1_v__reg[2]|Q_net ), .F1(\cal1_u54_XORCI_2|SUM_net ), .F2(dummy_abc_38_), .F3(dummy_abc_39_) );
      defparam ii0752.CONFIG_DATA = 16'h9999;
      defparam ii0752.PLACE_LOCATION = "NONE";
      defparam ii0752.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0753 ( .DX(nn0753), .F0(\cal1_v__reg[3]|Q_net ), .F1(\cal1_u54_XORCI_3|SUM_net ), .F2(dummy_abc_40_), .F3(dummy_abc_41_) );
      defparam ii0753.CONFIG_DATA = 16'h9999;
      defparam ii0753.PLACE_LOCATION = "NONE";
      defparam ii0753.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0754 ( .DX(nn0754), .F0(\cal1_v__reg[4]|Q_net ), .F1(\cal1_u54_XORCI_4|SUM_net ), .F2(dummy_abc_42_), .F3(dummy_abc_43_) );
      defparam ii0754.CONFIG_DATA = 16'h9999;
      defparam ii0754.PLACE_LOCATION = "NONE";
      defparam ii0754.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0755 ( .DX(nn0755), .F0(\cal1_v__reg[5]|Q_net ), .F1(\cal1_u54_XORCI_5|SUM_net ), .F2(dummy_abc_44_), .F3(dummy_abc_45_) );
      defparam ii0755.CONFIG_DATA = 16'h9999;
      defparam ii0755.PLACE_LOCATION = "NONE";
      defparam ii0755.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0756 ( .DX(nn0756), .F0(\cal1_u54_XORCI_6|SUM_net ), .F1(dummy_abc_46_), .F2(dummy_abc_47_), .F3(dummy_abc_48_) );
      defparam ii0756.CONFIG_DATA = 16'h5555;
      defparam ii0756.PLACE_LOCATION = "NONE";
      defparam ii0756.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7_5_ ( 
        .CA( {\cal1_u54_XORCI_6|SUM_net , \cal1_u54_XORCI_5|SUM_net , 
              \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_3|SUM_net , \cal1_u54_XORCI_2|SUM_net , 
              \cal1_u54_XORCI_1|SUM_net , \cal1_uPreF__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_885_ ), 
        .DX( {nn0756, nn0755, nn0754, nn0753, nn0752, nn0751, nn0750} ), 
        .SUM( {\cal1_u55_XORCI_6|SUM_net , \cal1_u55_XORCI_5|SUM_net , 
              \cal1_u55_XORCI_4|SUM_net , \cal1_u55_XORCI_3|SUM_net , \cal1_u55_XORCI_2|SUM_net , 
              \cal1_u55_XORCI_1|SUM_net , \cal1_u55_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0766 ( .DX(nn0766), .F0(\a_mac_out[7]_cal1_u134_mac ), .F1(\cal1_u55_XORCI_1|SUM_net ), .F2(dummy_abc_49_), .F3(dummy_abc_50_) );
      defparam ii0766.CONFIG_DATA = 16'h6666;
      defparam ii0766.PLACE_LOCATION = "NONE";
      defparam ii0766.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0767 ( .DX(nn0767), .F0(\a_mac_out[8]_cal1_u134_mac ), .F1(\cal1_u55_XORCI_2|SUM_net ), .F2(dummy_abc_51_), .F3(dummy_abc_52_) );
      defparam ii0767.CONFIG_DATA = 16'h6666;
      defparam ii0767.PLACE_LOCATION = "NONE";
      defparam ii0767.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0768 ( .DX(nn0768), .F0(\a_mac_out[9]_cal1_u134_mac ), .F1(\cal1_u55_XORCI_3|SUM_net ), .F2(dummy_abc_53_), .F3(dummy_abc_54_) );
      defparam ii0768.CONFIG_DATA = 16'h6666;
      defparam ii0768.PLACE_LOCATION = "NONE";
      defparam ii0768.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0769 ( .DX(nn0769), .F0(\a_mac_out[10]_cal1_u134_mac ), .F1(\cal1_u55_XORCI_4|SUM_net ), .F2(dummy_abc_55_), .F3(dummy_abc_56_) );
      defparam ii0769.CONFIG_DATA = 16'h6666;
      defparam ii0769.PLACE_LOCATION = "NONE";
      defparam ii0769.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0770 ( .DX(nn0770), .F0(\a_mac_out[11]_cal1_u134_mac ), .F1(\cal1_u55_XORCI_5|SUM_net ), .F2(dummy_abc_57_), .F3(dummy_abc_58_) );
      defparam ii0770.CONFIG_DATA = 16'h6666;
      defparam ii0770.PLACE_LOCATION = "NONE";
      defparam ii0770.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0771 ( .DX(nn0771), .F0(\cal1_u55_XORCI_6|SUM_net ), .F1(dummy_abc_59_), .F2(dummy_abc_60_), .F3(dummy_abc_61_) );
      defparam ii0771.CONFIG_DATA = 16'hAAAA;
      defparam ii0771.PLACE_LOCATION = "NONE";
      defparam ii0771.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7 ( 
        .CA( {a_acc_en_cal1_u134_mac, \a_mac_out[11]_cal1_u134_mac , 
              \a_mac_out[10]_cal1_u134_mac , \a_mac_out[9]_cal1_u134_mac , \a_mac_out[8]_cal1_u134_mac , 
              \a_mac_out[7]_cal1_u134_mac , \a_mac_out[6]_cal1_u134_mac } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_883_ ), 
        .DX( {nn0771, nn0770, nn0769, nn0768, nn0767, nn0766, nn0732} ), 
        .SUM( {\cal1_u133_XORCI_6|SUM_net , \cal1_u133_XORCI_5|SUM_net , 
              \cal1_u133_XORCI_4|SUM_net , \cal1_u133_XORCI_3|SUM_net , \cal1_u133_XORCI_2|SUM_net , 
              \cal1_u133_XORCI_1|SUM_net , \cal1_u133_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0781 ( .DX(\a_dinx[0]_cal1_u136_mac ), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[0]|Q_net ), .F2(dummy_abc_62_), .F3(dummy_abc_63_) );
      defparam ii0781.CONFIG_DATA = 16'h6666;
      defparam ii0781.PLACE_LOCATION = "NONE";
      defparam ii0781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0782 ( .DX(\a_dinx[0]_cal1_u137_mac ), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_abc_64_), .F3(dummy_abc_65_) );
      defparam ii0782.CONFIG_DATA = 16'h6666;
      defparam ii0782.PLACE_LOCATION = "NONE";
      defparam ii0782.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0783 ( .DX(\a_dinx[1]_cal1_u136_mac ), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\a_mac_out[7]_cal1_u134_mac ), .F2(\cal1_uPreF__reg[0]|Q_net ), .F3(\cal1_uPreF__reg[1]|Q_net ) );
      defparam ii0783.CONFIG_DATA = 16'h39C6;
      defparam ii0783.PLACE_LOCATION = "NONE";
      defparam ii0783.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0784 ( .DX(\a_dinx[1]_cal1_u137_mac ), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\a_mac_out[7]_cal1_u134_mac ), .F2(\cal1_v__reg[0]|Q_net ), .F3(\cal1_v__reg[1]|Q_net ) );
      defparam ii0784.CONFIG_DATA = 16'h39C6;
      defparam ii0784.PLACE_LOCATION = "NONE";
      defparam ii0784.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0785 ( .DX(nn0785), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\a_mac_out[7]_cal1_u134_mac ), .F2(\cal1_uPreF__reg[0]|Q_net ), .F3(\cal1_uPreF__reg[1]|Q_net ) );
      defparam ii0785.CONFIG_DATA = 16'h08CE;
      defparam ii0785.PLACE_LOCATION = "NONE";
      defparam ii0785.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0786 ( .DX(\a_dinx[2]_cal1_u136_mac ), .F0(\a_mac_out[8]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[2]|Q_net ), .F2(nn0785), .F3(dummy_abc_66_) );
      defparam ii0786.CONFIG_DATA = 16'h9696;
      defparam ii0786.PLACE_LOCATION = "NONE";
      defparam ii0786.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0787 ( .DX(nn0787), .F0(\a_mac_out[6]_cal1_u134_mac ), .F1(\a_mac_out[7]_cal1_u134_mac ), .F2(\cal1_v__reg[0]|Q_net ), .F3(\cal1_v__reg[1]|Q_net ) );
      defparam ii0787.CONFIG_DATA = 16'h08CE;
      defparam ii0787.PLACE_LOCATION = "NONE";
      defparam ii0787.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0788 ( .DX(\a_dinx[2]_cal1_u137_mac ), .F0(\a_mac_out[8]_cal1_u134_mac ), .F1(\cal1_v__reg[2]|Q_net ), .F2(nn0787), .F3(dummy_abc_67_) );
      defparam ii0788.CONFIG_DATA = 16'h9696;
      defparam ii0788.PLACE_LOCATION = "NONE";
      defparam ii0788.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0789 ( .DX(nn0789), .F0(\a_mac_out[8]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[2]|Q_net ), .F2(nn0785), .F3(dummy_abc_68_) );
      defparam ii0789.CONFIG_DATA = 16'h4D4D;
      defparam ii0789.PLACE_LOCATION = "NONE";
      defparam ii0789.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0790 ( .DX(\a_dinx[3]_cal1_u136_mac ), .F0(\a_mac_out[9]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[3]|Q_net ), .F2(nn0789), .F3(dummy_abc_69_) );
      defparam ii0790.CONFIG_DATA = 16'h6969;
      defparam ii0790.PLACE_LOCATION = "NONE";
      defparam ii0790.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0791 ( .DX(nn0791), .F0(\a_mac_out[8]_cal1_u134_mac ), .F1(\cal1_v__reg[2]|Q_net ), .F2(nn0787), .F3(dummy_abc_70_) );
      defparam ii0791.CONFIG_DATA = 16'h4D4D;
      defparam ii0791.PLACE_LOCATION = "NONE";
      defparam ii0791.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0792 ( .DX(\a_dinx[3]_cal1_u137_mac ), .F0(\a_mac_out[9]_cal1_u134_mac ), .F1(\cal1_v__reg[3]|Q_net ), .F2(nn0791), .F3(dummy_abc_71_) );
      defparam ii0792.CONFIG_DATA = 16'h6969;
      defparam ii0792.PLACE_LOCATION = "NONE";
      defparam ii0792.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0793 ( .DX(nn0793), .F0(\a_mac_out[9]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[3]|Q_net ), .F2(nn0789), .F3(dummy_abc_72_) );
      defparam ii0793.CONFIG_DATA = 16'h2B2B;
      defparam ii0793.PLACE_LOCATION = "NONE";
      defparam ii0793.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0794 ( .DX(\a_dinx[4]_cal1_u136_mac ), .F0(\a_mac_out[10]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[4]|Q_net ), .F2(nn0793), .F3(dummy_abc_73_) );
      defparam ii0794.CONFIG_DATA = 16'h9696;
      defparam ii0794.PLACE_LOCATION = "NONE";
      defparam ii0794.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0795 ( .DX(nn0795), .F0(\a_mac_out[9]_cal1_u134_mac ), .F1(\cal1_v__reg[3]|Q_net ), .F2(nn0791), .F3(dummy_abc_74_) );
      defparam ii0795.CONFIG_DATA = 16'h2B2B;
      defparam ii0795.PLACE_LOCATION = "NONE";
      defparam ii0795.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0796 ( .DX(\a_dinx[4]_cal1_u137_mac ), .F0(\a_mac_out[10]_cal1_u134_mac ), .F1(\cal1_v__reg[4]|Q_net ), .F2(nn0795), .F3(dummy_abc_75_) );
      defparam ii0796.CONFIG_DATA = 16'h9696;
      defparam ii0796.PLACE_LOCATION = "NONE";
      defparam ii0796.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0797 ( .DX(nn0797), .F0(\a_mac_out[11]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[5]|Q_net ), .F2(dummy_abc_76_), .F3(dummy_abc_77_) );
      defparam ii0797.CONFIG_DATA = 16'h6666;
      defparam ii0797.PLACE_LOCATION = "NONE";
      defparam ii0797.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0798 ( .DX(\a_dinx[5]_cal1_u136_mac ), .F0(\a_mac_out[10]_cal1_u134_mac ), .F1(\cal1_uPreF__reg[4]|Q_net ), .F2(nn0793), .F3(nn0797) );
      defparam ii0798.CONFIG_DATA = 16'h4DB2;
      defparam ii0798.PLACE_LOCATION = "NONE";
      defparam ii0798.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0799 ( .DX(nn0799), .F0(\a_mac_out[11]_cal1_u134_mac ), .F1(\cal1_v__reg[5]|Q_net ), .F2(dummy_abc_78_), .F3(dummy_abc_79_) );
      defparam ii0799.CONFIG_DATA = 16'h6666;
      defparam ii0799.PLACE_LOCATION = "NONE";
      defparam ii0799.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0800 ( .DX(\a_dinx[5]_cal1_u137_mac ), .F0(\a_mac_out[10]_cal1_u134_mac ), .F1(\cal1_v__reg[4]|Q_net ), .F2(nn0795), .F3(nn0799) );
      defparam ii0800.CONFIG_DATA = 16'h4DB2;
      defparam ii0800.PLACE_LOCATION = "NONE";
      defparam ii0800.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0801 ( .DX(nn0801), .F0(\cal1_enforceJmp__reg|Q_net ), .F1(\cal1_jmp1Normal__reg|Q_net ), .F2(dummy_abc_80_), .F3(dummy_abc_81_) );
      defparam ii0801.CONFIG_DATA = 16'h1111;
      defparam ii0801.PLACE_LOCATION = "NONE";
      defparam ii0801.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0802 ( .DX(nn0802), .F0(rst), .F1(u4168_or2_41__I0), .F2(u4168_or2_41__I0_5_), .F3(nn0801) );
      defparam ii0802.CONFIG_DATA = 16'h1105;
      defparam ii0802.PLACE_LOCATION = "NONE";
      defparam ii0802.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0803 ( .DX(nn0803), .F0(rst), .F1(\cal1_jmp2Normal__reg|Q_net ), .F2(nn0801), .F3(nn0802) );
      defparam ii0803.CONFIG_DATA = 16'h00BA;
      defparam ii0803.PLACE_LOCATION = "NONE";
      defparam ii0803.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0804 ( .DX(nn0804), .F0(\c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_82_) );
      defparam ii0804.CONFIG_DATA = 16'hCACA;
      defparam ii0804.PLACE_LOCATION = "NONE";
      defparam ii0804.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0805 ( .DX(nn0805), .F0(u4168_or2_41__I0_5_), .F1(u4168_or2_41__IN), .F2(\cal1_jmp2Normal__reg|Q_net ), .F3(nn0801) );
      defparam ii0805.CONFIG_DATA = 16'hC0AA;
      defparam ii0805.PLACE_LOCATION = "NONE";
      defparam ii0805.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0806 ( .DX(nn0806), .F0(u4168_or2_41__IN), .F1(nn0802), .F2(nn0805), .F3(dummy_abc_83_) );
      defparam ii0806.CONFIG_DATA = 16'h0808;
      defparam ii0806.PLACE_LOCATION = "NONE";
      defparam ii0806.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0807 ( .DX(nn0807), .F0(\c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0807.CONFIG_DATA = 16'h35FF;
      defparam ii0807.PLACE_LOCATION = "NONE";
      defparam ii0807.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0808 ( .DX(\a_diny[0]_cal1_u135_mac ), .F0(nn0803), .F1(nn0804), .F2(nn0807), .F3(dummy_abc_84_) );
      defparam ii0808.CONFIG_DATA = 16'h8F8F;
      defparam ii0808.PLACE_LOCATION = "NONE";
      defparam ii0808.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0809 ( .DX(nn0809), .F0(\c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_85_) );
      defparam ii0809.CONFIG_DATA = 16'h3535;
      defparam ii0809.PLACE_LOCATION = "NONE";
      defparam ii0809.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0810 ( .DX(nn0810), .F0(\c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0810.CONFIG_DATA = 16'h35FF;
      defparam ii0810.PLACE_LOCATION = "NONE";
      defparam ii0810.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0811 ( .DX(\a_diny[0]_cal1_u136_mac ), .F0(nn0803), .F1(nn0809), .F2(nn0810), .F3(dummy_abc_86_) );
      defparam ii0811.CONFIG_DATA = 16'h2F2F;
      defparam ii0811.PLACE_LOCATION = "NONE";
      defparam ii0811.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0812 ( .DX(nn0812), .F0(xBgn[0]), .F1(xEnd[0]), .F2(dummy_abc_87_), .F3(dummy_abc_88_) );
      defparam ii0812.CONFIG_DATA = 16'h6666;
      defparam ii0812.PLACE_LOCATION = "NONE";
      defparam ii0812.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0813 ( .DX(nn0813), .F0(\cal1_v__reg[6]|Q_net ), .F1(nn0812), .F2(dummy_abc_89_), .F3(dummy_abc_90_) );
      defparam ii0813.CONFIG_DATA = 16'h6666;
      defparam ii0813.PLACE_LOCATION = "NONE";
      defparam ii0813.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0814 ( .DX(nn0814), .F0(nn0812), .F1(dummy_abc_91_), .F2(dummy_abc_92_), .F3(dummy_abc_93_) );
      defparam ii0814.CONFIG_DATA = 16'h5555;
      defparam ii0814.PLACE_LOCATION = "NONE";
      defparam ii0814.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0815 ( .DX(nn0815), .F0(xBgn[1]), .F1(xEnd[1]), .F2(dummy_abc_94_), .F3(dummy_abc_95_) );
      defparam ii0815.CONFIG_DATA = 16'h9999;
      defparam ii0815.PLACE_LOCATION = "NONE";
      defparam ii0815.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0816 ( .DX(nn0816), .F0(xBgn[2]), .F1(xEnd[2]), .F2(dummy_abc_96_), .F3(dummy_abc_97_) );
      defparam ii0816.CONFIG_DATA = 16'h9999;
      defparam ii0816.PLACE_LOCATION = "NONE";
      defparam ii0816.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0817 ( .DX(nn0817), .F0(xBgn[3]), .F1(xEnd[3]), .F2(dummy_abc_98_), .F3(dummy_abc_99_) );
      defparam ii0817.CONFIG_DATA = 16'h9999;
      defparam ii0817.PLACE_LOCATION = "NONE";
      defparam ii0817.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0818 ( .DX(nn0818), .F0(xBgn[4]), .F1(xEnd[4]), .F2(dummy_abc_100_), .F3(dummy_abc_101_) );
      defparam ii0818.CONFIG_DATA = 16'h9999;
      defparam ii0818.PLACE_LOCATION = "NONE";
      defparam ii0818.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0819 ( .DX(nn0819), .F0(xBgn[5]), .F1(xEnd[5]), .F2(dummy_abc_102_), .F3(dummy_abc_103_) );
      defparam ii0819.CONFIG_DATA = 16'h9999;
      defparam ii0819.PLACE_LOCATION = "NONE";
      defparam ii0819.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0820 ( .DX(nn0820), .F0(xBgn[6]), .F1(xEnd[6]), .F2(dummy_abc_104_), .F3(dummy_abc_105_) );
      defparam ii0820.CONFIG_DATA = 16'h9999;
      defparam ii0820.PLACE_LOCATION = "NONE";
      defparam ii0820.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0821 ( .DX(nn0821), .F0(xBgn[7]), .F1(xEnd[7]), .F2(dummy_abc_106_), .F3(dummy_abc_107_) );
      defparam ii0821.CONFIG_DATA = 16'h9999;
      defparam ii0821.PLACE_LOCATION = "NONE";
      defparam ii0821.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0822 ( .DX(nn0822), .F0(xBgn[8]), .F1(xEnd[8]), .F2(dummy_abc_108_), .F3(dummy_abc_109_) );
      defparam ii0822.CONFIG_DATA = 16'h9999;
      defparam ii0822.PLACE_LOCATION = "NONE";
      defparam ii0822.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0823 ( .DX(nn0823), .F0(xBgn[9]), .F1(xEnd[9]), .F2(dummy_abc_110_), .F3(dummy_abc_111_) );
      defparam ii0823.CONFIG_DATA = 16'h9999;
      defparam ii0823.PLACE_LOCATION = "NONE";
      defparam ii0823.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0824 ( .DX(nn0824), .F0(xBgn[10]), .F1(xEnd[10]), .F2(dummy_abc_112_), .F3(dummy_abc_113_) );
      defparam ii0824.CONFIG_DATA = 16'h9999;
      defparam ii0824.PLACE_LOCATION = "NONE";
      defparam ii0824.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0825 ( .DX(nn0825), .F0(dummy_abc_114_), .F1(dummy_abc_115_), .F2(dummy_abc_116_), .F3(dummy_abc_117_) );
      defparam ii0825.CONFIG_DATA = 16'hFFFF;
      defparam ii0825.PLACE_LOCATION = "NONE";
      defparam ii0825.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_88_ ( 
        .CA( {a_acc_en_cal1_u134_mac, xEnd[10], xEnd[9], xEnd[8], xEnd[7], 
              xEnd[6], xEnd[5], xEnd[4], xEnd[3], xEnd[2], xEnd[1], xEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_119_ ), 
        .DX( {nn0825, nn0824, nn0823, nn0822, nn0821, nn0820, nn0819, nn0818, 
              nn0817, nn0816, nn0815, nn0814} ), 
        .SUM( {\u2_XORCI_11|SUM_net , \u2_XORCI_10|SUM_net , \u2_XORCI_9|SUM_net , 
              \u2_XORCI_8|SUM_net , \u2_XORCI_7|SUM_net , \u2_XORCI_6|SUM_net , 
              \u2_XORCI_5|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_3|SUM_net , 
              \u2_XORCI_2|SUM_net , \u2_XORCI_1|SUM_net , \u2_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0840 ( .DX(nn0840), .F0(xBgn[0]), .F1(xEnd[0]), .F2(dummy_abc_118_), .F3(dummy_abc_119_) );
      defparam ii0840.CONFIG_DATA = 16'h6666;
      defparam ii0840.PLACE_LOCATION = "NONE";
      defparam ii0840.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0841 ( .DX(nn0841), .F0(\u2_XORCI_1|SUM_net ), .F1(dummy_abc_120_), .F2(dummy_abc_121_), .F3(dummy_abc_122_) );
      defparam ii0841.CONFIG_DATA = 16'h5555;
      defparam ii0841.PLACE_LOCATION = "NONE";
      defparam ii0841.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0842 ( .DX(nn0842), .F0(\u2_XORCI_2|SUM_net ), .F1(dummy_abc_123_), .F2(dummy_abc_124_), .F3(dummy_abc_125_) );
      defparam ii0842.CONFIG_DATA = 16'h5555;
      defparam ii0842.PLACE_LOCATION = "NONE";
      defparam ii0842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0843 ( .DX(nn0843), .F0(\u2_XORCI_3|SUM_net ), .F1(dummy_abc_126_), .F2(dummy_abc_127_), .F3(dummy_abc_128_) );
      defparam ii0843.CONFIG_DATA = 16'h5555;
      defparam ii0843.PLACE_LOCATION = "NONE";
      defparam ii0843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0844 ( .DX(nn0844), .F0(\u2_XORCI_4|SUM_net ), .F1(dummy_abc_129_), .F2(dummy_abc_130_), .F3(dummy_abc_131_) );
      defparam ii0844.CONFIG_DATA = 16'h5555;
      defparam ii0844.PLACE_LOCATION = "NONE";
      defparam ii0844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0845 ( .DX(nn0845), .F0(\u2_XORCI_5|SUM_net ), .F1(dummy_abc_132_), .F2(dummy_abc_133_), .F3(dummy_abc_134_) );
      defparam ii0845.CONFIG_DATA = 16'h5555;
      defparam ii0845.PLACE_LOCATION = "NONE";
      defparam ii0845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0846 ( .DX(nn0846), .F0(\u2_XORCI_6|SUM_net ), .F1(dummy_abc_135_), .F2(dummy_abc_136_), .F3(dummy_abc_137_) );
      defparam ii0846.CONFIG_DATA = 16'h5555;
      defparam ii0846.PLACE_LOCATION = "NONE";
      defparam ii0846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0847 ( .DX(nn0847), .F0(\u2_XORCI_7|SUM_net ), .F1(dummy_abc_138_), .F2(dummy_abc_139_), .F3(dummy_abc_140_) );
      defparam ii0847.CONFIG_DATA = 16'h5555;
      defparam ii0847.PLACE_LOCATION = "NONE";
      defparam ii0847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0848 ( .DX(nn0848), .F0(\u2_XORCI_8|SUM_net ), .F1(dummy_abc_141_), .F2(dummy_abc_142_), .F3(dummy_abc_143_) );
      defparam ii0848.CONFIG_DATA = 16'h5555;
      defparam ii0848.PLACE_LOCATION = "NONE";
      defparam ii0848.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0849 ( .DX(nn0849), .F0(\u2_XORCI_9|SUM_net ), .F1(dummy_abc_144_), .F2(dummy_abc_145_), .F3(dummy_abc_146_) );
      defparam ii0849.CONFIG_DATA = 16'h5555;
      defparam ii0849.PLACE_LOCATION = "NONE";
      defparam ii0849.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0850 ( .DX(nn0850), .F0(\u2_XORCI_10|SUM_net ), .F1(dummy_abc_147_), .F2(dummy_abc_148_), .F3(dummy_abc_149_) );
      defparam ii0850.CONFIG_DATA = 16'h5555;
      defparam ii0850.PLACE_LOCATION = "NONE";
      defparam ii0850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0851 ( .DX(nn0851), .F0(dummy_abc_150_), .F1(dummy_abc_151_), .F2(dummy_abc_152_), .F3(dummy_abc_153_) );
      defparam ii0851.CONFIG_DATA = 16'h0000;
      defparam ii0851.PLACE_LOCATION = "NONE";
      defparam ii0851.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_89_ ( 
        .CA( {\u2_XORCI_11|SUM_net , \u2_XORCI_10|SUM_net , \u2_XORCI_9|SUM_net , 
              \u2_XORCI_8|SUM_net , \u2_XORCI_7|SUM_net , \u2_XORCI_6|SUM_net , 
              \u2_XORCI_5|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_3|SUM_net , 
              \u2_XORCI_2|SUM_net , \u2_XORCI_1|SUM_net , nn0812} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_120_ ), 
        .DX( {nn0851, nn0850, nn0849, nn0848, nn0847, nn0846, nn0845, nn0844, 
              nn0843, nn0842, nn0841, nn0840} ), 
        .SUM( {dummy_121_, \u3_XORCI_10|SUM_net , \u3_XORCI_9|SUM_net , 
              \u3_XORCI_8|SUM_net , \u3_XORCI_7|SUM_net , \u3_XORCI_6|SUM_net , 
              \u3_XORCI_5|SUM_net , \u3_XORCI_4|SUM_net , \u3_XORCI_3|SUM_net , 
              \u3_XORCI_2|SUM_net , \u3_XORCI_1|SUM_net , \u3_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0866 ( .DX(nn0866), .F0(\cal1_v__reg[7]|Q_net ), .F1(\u3_XORCI_1|SUM_net ), .F2(dummy_abc_154_), .F3(dummy_abc_155_) );
      defparam ii0866.CONFIG_DATA = 16'h9999;
      defparam ii0866.PLACE_LOCATION = "NONE";
      defparam ii0866.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0867 ( .DX(nn0867), .F0(\cal1_v__reg[8]|Q_net ), .F1(\u3_XORCI_2|SUM_net ), .F2(dummy_abc_156_), .F3(dummy_abc_157_) );
      defparam ii0867.CONFIG_DATA = 16'h9999;
      defparam ii0867.PLACE_LOCATION = "NONE";
      defparam ii0867.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0868 ( .DX(nn0868), .F0(\cal1_v__reg[9]|Q_net ), .F1(\u3_XORCI_3|SUM_net ), .F2(dummy_abc_158_), .F3(dummy_abc_159_) );
      defparam ii0868.CONFIG_DATA = 16'h9999;
      defparam ii0868.PLACE_LOCATION = "NONE";
      defparam ii0868.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0869 ( .DX(nn0869), .F0(\cal1_v__reg[10]|Q_net ), .F1(\u3_XORCI_4|SUM_net ), .F2(dummy_abc_160_), .F3(dummy_abc_161_) );
      defparam ii0869.CONFIG_DATA = 16'h9999;
      defparam ii0869.PLACE_LOCATION = "NONE";
      defparam ii0869.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0870 ( .DX(nn0870), .F0(\cal1_v__reg[11]|Q_net ), .F1(\u3_XORCI_5|SUM_net ), .F2(dummy_abc_162_), .F3(dummy_abc_163_) );
      defparam ii0870.CONFIG_DATA = 16'h9999;
      defparam ii0870.PLACE_LOCATION = "NONE";
      defparam ii0870.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0871 ( .DX(nn0871), .F0(\cal1_v__reg[12]|Q_net ), .F1(\u3_XORCI_6|SUM_net ), .F2(dummy_abc_164_), .F3(dummy_abc_165_) );
      defparam ii0871.CONFIG_DATA = 16'h9999;
      defparam ii0871.PLACE_LOCATION = "NONE";
      defparam ii0871.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0872 ( .DX(nn0872), .F0(\cal1_v__reg[13]|Q_net ), .F1(\u3_XORCI_7|SUM_net ), .F2(dummy_abc_166_), .F3(dummy_abc_167_) );
      defparam ii0872.CONFIG_DATA = 16'h9999;
      defparam ii0872.PLACE_LOCATION = "NONE";
      defparam ii0872.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0873 ( .DX(nn0873), .F0(\cal1_v__reg[14]|Q_net ), .F1(\u3_XORCI_8|SUM_net ), .F2(dummy_abc_168_), .F3(dummy_abc_169_) );
      defparam ii0873.CONFIG_DATA = 16'h9999;
      defparam ii0873.PLACE_LOCATION = "NONE";
      defparam ii0873.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0874 ( .DX(nn0874), .F0(\cal1_v__reg[15]|Q_net ), .F1(\u3_XORCI_9|SUM_net ), .F2(dummy_abc_170_), .F3(dummy_abc_171_) );
      defparam ii0874.CONFIG_DATA = 16'h9999;
      defparam ii0874.PLACE_LOCATION = "NONE";
      defparam ii0874.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0875 ( .DX(nn0875), .F0(\cal1_v__reg[16]|Q_net ), .F1(\u3_XORCI_10|SUM_net ), .F2(dummy_abc_172_), .F3(dummy_abc_173_) );
      defparam ii0875.CONFIG_DATA = 16'h9999;
      defparam ii0875.PLACE_LOCATION = "NONE";
      defparam ii0875.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0876 ( .DX(nn0876), .F0(dummy_abc_174_), .F1(dummy_abc_175_), .F2(dummy_abc_176_), .F3(dummy_abc_177_) );
      defparam ii0876.CONFIG_DATA = 16'hFFFF;
      defparam ii0876.PLACE_LOCATION = "NONE";
      defparam ii0876.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_8_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \cal1_v__reg[16]|Q_net , 
              \cal1_v__reg[15]|Q_net , \cal1_v__reg[14]|Q_net , \cal1_v__reg[13]|Q_net , 
              \cal1_v__reg[12]|Q_net , \cal1_v__reg[11]|Q_net , \cal1_v__reg[10]|Q_net , 
              \cal1_v__reg[9]|Q_net , \cal1_v__reg[8]|Q_net , \cal1_v__reg[7]|Q_net , 
              \cal1_v__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_123_ ), 
        .DX( {nn0876, nn0875, nn0874, nn0873, nn0872, nn0871, nn0870, nn0869, 
              nn0868, nn0867, nn0866, nn0813} ), 
        .SUM( {\cal1_u63_XORCI_11|SUM_net , dummy_124_, dummy_125_, dummy_126_, 
              dummy_127_, dummy_128_, dummy_129_, dummy_130_, dummy_131_, dummy_132_, 
              dummy_133_, dummy_134_} )
      );
    CS_LUT4_PRIM ii0891 ( .DX(nn0891), .F0(\fifo1_ram_inst_1_aa_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0803), .F3(dummy_abc_178_) );
      defparam ii0891.CONFIG_DATA = 16'h1010;
      defparam ii0891.PLACE_LOCATION = "NONE";
      defparam ii0891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0892 ( .DX(nn0892), .F0(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0806), .F3(dummy_abc_179_) );
      defparam ii0892.CONFIG_DATA = 16'h1010;
      defparam ii0892.PLACE_LOCATION = "NONE";
      defparam ii0892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0893 ( .DX(nn0893), .F0(\fifo1_ram_inst_1_aa_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0803), .F3(dummy_abc_180_) );
      defparam ii0893.CONFIG_DATA = 16'h2020;
      defparam ii0893.PLACE_LOCATION = "NONE";
      defparam ii0893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0894 ( .DX(nn0894), .F0(\c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0892), .F3(nn0893) );
      defparam ii0894.CONFIG_DATA = 16'h135F;
      defparam ii0894.PLACE_LOCATION = "NONE";
      defparam ii0894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0895 ( .DX(nn0895), .F0(\c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0891), .F2(nn0894), .F3(dummy_abc_181_) );
      defparam ii0895.CONFIG_DATA = 16'h7070;
      defparam ii0895.PLACE_LOCATION = "NONE";
      defparam ii0895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0896 ( .DX(\a_diny[0]_cal1_u137_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u135_mac ), .F2(nn0895), .F3(dummy_abc_182_) );
      defparam ii0896.CONFIG_DATA = 16'h8F8F;
      defparam ii0896.PLACE_LOCATION = "NONE";
      defparam ii0896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0897 ( .DX(nn0897), .F0(\fifo1_ram_inst_1_ab_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0803), .F3(dummy_abc_183_) );
      defparam ii0897.CONFIG_DATA = 16'h2020;
      defparam ii0897.PLACE_LOCATION = "NONE";
      defparam ii0897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0898 ( .DX(nn0898), .F0(\fifo1_ram_inst_1_ab_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0803), .F3(dummy_abc_184_) );
      defparam ii0898.CONFIG_DATA = 16'h1010;
      defparam ii0898.PLACE_LOCATION = "NONE";
      defparam ii0898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0899 ( .DX(nn0899), .F0(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F1(dummy_123_), .F2(nn0806), .F3(dummy_abc_185_) );
      defparam ii0899.CONFIG_DATA = 16'h1010;
      defparam ii0899.PLACE_LOCATION = "NONE";
      defparam ii0899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0900 ( .DX(nn0900), .F0(\c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0898), .F3(nn0899) );
      defparam ii0900.CONFIG_DATA = 16'h153F;
      defparam ii0900.PLACE_LOCATION = "NONE";
      defparam ii0900.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0901 ( .DX(nn0901), .F0(\c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0897), .F2(nn0900), .F3(dummy_abc_186_) );
      defparam ii0901.CONFIG_DATA = 16'h7070;
      defparam ii0901.PLACE_LOCATION = "NONE";
      defparam ii0901.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0902 ( .DX(\a_diny[0]_cal1_u138_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u136_mac ), .F2(nn0901), .F3(dummy_abc_187_) );
      defparam ii0902.CONFIG_DATA = 16'h8F8F;
      defparam ii0902.PLACE_LOCATION = "NONE";
      defparam ii0902.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0903 ( .DX(nn0903), .F0(\c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_188_) );
      defparam ii0903.CONFIG_DATA = 16'hCACA;
      defparam ii0903.PLACE_LOCATION = "NONE";
      defparam ii0903.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0904 ( .DX(nn0904), .F0(\c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0904.CONFIG_DATA = 16'h35FF;
      defparam ii0904.PLACE_LOCATION = "NONE";
      defparam ii0904.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0905 ( .DX(\a_diny[0]_cal1_u139_mac ), .F0(nn0803), .F1(nn0903), .F2(nn0904), .F3(dummy_abc_189_) );
      defparam ii0905.CONFIG_DATA = 16'h8F8F;
      defparam ii0905.PLACE_LOCATION = "NONE";
      defparam ii0905.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0906 ( .DX(nn0906), .F0(\c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_190_) );
      defparam ii0906.CONFIG_DATA = 16'h3535;
      defparam ii0906.PLACE_LOCATION = "NONE";
      defparam ii0906.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0907 ( .DX(nn0907), .F0(\c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0907.CONFIG_DATA = 16'h35FF;
      defparam ii0907.PLACE_LOCATION = "NONE";
      defparam ii0907.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0908 ( .DX(\a_diny[0]_cal1_u140_mac ), .F0(nn0803), .F1(nn0906), .F2(nn0907), .F3(dummy_abc_191_) );
      defparam ii0908.CONFIG_DATA = 16'h2F2F;
      defparam ii0908.PLACE_LOCATION = "NONE";
      defparam ii0908.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0909 ( .DX(nn0909), .F0(\c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0891) );
      defparam ii0909.CONFIG_DATA = 16'h135F;
      defparam ii0909.PLACE_LOCATION = "NONE";
      defparam ii0909.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0910 ( .DX(nn0910), .F0(\c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0893), .F2(nn0909), .F3(dummy_abc_192_) );
      defparam ii0910.CONFIG_DATA = 16'h7070;
      defparam ii0910.PLACE_LOCATION = "NONE";
      defparam ii0910.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0911 ( .DX(\a_diny[0]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u139_mac ), .F2(nn0910), .F3(dummy_abc_193_) );
      defparam ii0911.CONFIG_DATA = 16'h8F8F;
      defparam ii0911.PLACE_LOCATION = "NONE";
      defparam ii0911.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0912 ( .DX(nn0912), .F0(\c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0899) );
      defparam ii0912.CONFIG_DATA = 16'h153F;
      defparam ii0912.PLACE_LOCATION = "NONE";
      defparam ii0912.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0913 ( .DX(nn0913), .F0(\c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0897), .F2(nn0912), .F3(dummy_abc_194_) );
      defparam ii0913.CONFIG_DATA = 16'h7070;
      defparam ii0913.PLACE_LOCATION = "NONE";
      defparam ii0913.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0914 ( .DX(\a_diny[0]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u140_mac ), .F2(nn0913), .F3(dummy_abc_195_) );
      defparam ii0914.CONFIG_DATA = 16'h8F8F;
      defparam ii0914.PLACE_LOCATION = "NONE";
      defparam ii0914.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0915 ( .DX(nn0915), .F0(\c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_196_) );
      defparam ii0915.CONFIG_DATA = 16'h3535;
      defparam ii0915.PLACE_LOCATION = "NONE";
      defparam ii0915.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0916 ( .DX(nn0916), .F0(\c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0916.CONFIG_DATA = 16'h35FF;
      defparam ii0916.PLACE_LOCATION = "NONE";
      defparam ii0916.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0917 ( .DX(\a_diny[0]_cal1_u143_mac ), .F0(nn0803), .F1(nn0915), .F2(nn0916), .F3(dummy_abc_197_) );
      defparam ii0917.CONFIG_DATA = 16'h2F2F;
      defparam ii0917.PLACE_LOCATION = "NONE";
      defparam ii0917.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0918 ( .DX(nn0918), .F0(\c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_198_) );
      defparam ii0918.CONFIG_DATA = 16'hCACA;
      defparam ii0918.PLACE_LOCATION = "NONE";
      defparam ii0918.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0919 ( .DX(nn0919), .F0(\c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0919.CONFIG_DATA = 16'h35FF;
      defparam ii0919.PLACE_LOCATION = "NONE";
      defparam ii0919.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0920 ( .DX(\a_diny[0]_cal1_u144_mac ), .F0(nn0803), .F1(nn0918), .F2(nn0919), .F3(dummy_abc_199_) );
      defparam ii0920.CONFIG_DATA = 16'h8F8F;
      defparam ii0920.PLACE_LOCATION = "NONE";
      defparam ii0920.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0921 ( .DX(nn0921), .F0(\c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0893) );
      defparam ii0921.CONFIG_DATA = 16'h135F;
      defparam ii0921.PLACE_LOCATION = "NONE";
      defparam ii0921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0922 ( .DX(nn0922), .F0(\c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0891), .F2(nn0921), .F3(dummy_abc_200_) );
      defparam ii0922.CONFIG_DATA = 16'h7070;
      defparam ii0922.PLACE_LOCATION = "NONE";
      defparam ii0922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0923 ( .DX(\a_diny[0]_cal1_u145_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u143_mac ), .F2(nn0922), .F3(dummy_abc_201_) );
      defparam ii0923.CONFIG_DATA = 16'h8F8F;
      defparam ii0923.PLACE_LOCATION = "NONE";
      defparam ii0923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0924 ( .DX(nn0924), .F0(\c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0899) );
      defparam ii0924.CONFIG_DATA = 16'h153F;
      defparam ii0924.PLACE_LOCATION = "NONE";
      defparam ii0924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0925 ( .DX(nn0925), .F0(\c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0897), .F2(nn0924), .F3(dummy_abc_202_) );
      defparam ii0925.CONFIG_DATA = 16'h7070;
      defparam ii0925.PLACE_LOCATION = "NONE";
      defparam ii0925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0926 ( .DX(\a_diny[0]_cal1_u146_mac ), .F0(dummy_123_), .F1(\a_diny[0]_cal1_u144_mac ), .F2(nn0925), .F3(dummy_abc_203_) );
      defparam ii0926.CONFIG_DATA = 16'h8F8F;
      defparam ii0926.PLACE_LOCATION = "NONE";
      defparam ii0926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0927 ( .DX(nn0927), .F0(\c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_204_) );
      defparam ii0927.CONFIG_DATA = 16'h3535;
      defparam ii0927.PLACE_LOCATION = "NONE";
      defparam ii0927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0928 ( .DX(nn0928), .F0(\c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0928.CONFIG_DATA = 16'h35FF;
      defparam ii0928.PLACE_LOCATION = "NONE";
      defparam ii0928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0929 ( .DX(\a_diny[1]_cal1_u135_mac ), .F0(nn0803), .F1(nn0927), .F2(nn0928), .F3(dummy_abc_205_) );
      defparam ii0929.CONFIG_DATA = 16'h2F2F;
      defparam ii0929.PLACE_LOCATION = "NONE";
      defparam ii0929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0930 ( .DX(nn0930), .F0(\c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_206_) );
      defparam ii0930.CONFIG_DATA = 16'hCACA;
      defparam ii0930.PLACE_LOCATION = "NONE";
      defparam ii0930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0931 ( .DX(nn0931), .F0(\c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0931.CONFIG_DATA = 16'h35FF;
      defparam ii0931.PLACE_LOCATION = "NONE";
      defparam ii0931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0932 ( .DX(\a_diny[1]_cal1_u136_mac ), .F0(nn0803), .F1(nn0930), .F2(nn0931), .F3(dummy_abc_207_) );
      defparam ii0932.CONFIG_DATA = 16'h8F8F;
      defparam ii0932.PLACE_LOCATION = "NONE";
      defparam ii0932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0933 ( .DX(nn0933), .F0(\c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0891) );
      defparam ii0933.CONFIG_DATA = 16'h135F;
      defparam ii0933.PLACE_LOCATION = "NONE";
      defparam ii0933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0934 ( .DX(nn0934), .F0(\c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0893), .F2(nn0933), .F3(dummy_abc_208_) );
      defparam ii0934.CONFIG_DATA = 16'h7070;
      defparam ii0934.PLACE_LOCATION = "NONE";
      defparam ii0934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0935 ( .DX(\a_diny[1]_cal1_u137_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u135_mac ), .F2(nn0934), .F3(dummy_abc_209_) );
      defparam ii0935.CONFIG_DATA = 16'h8F8F;
      defparam ii0935.PLACE_LOCATION = "NONE";
      defparam ii0935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0936 ( .DX(nn0936), .F0(\c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0899) );
      defparam ii0936.CONFIG_DATA = 16'h153F;
      defparam ii0936.PLACE_LOCATION = "NONE";
      defparam ii0936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0937 ( .DX(nn0937), .F0(\c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0897), .F2(nn0936), .F3(dummy_abc_210_) );
      defparam ii0937.CONFIG_DATA = 16'h7070;
      defparam ii0937.PLACE_LOCATION = "NONE";
      defparam ii0937.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0938 ( .DX(\a_diny[1]_cal1_u138_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u136_mac ), .F2(nn0937), .F3(dummy_abc_211_) );
      defparam ii0938.CONFIG_DATA = 16'h8F8F;
      defparam ii0938.PLACE_LOCATION = "NONE";
      defparam ii0938.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0939 ( .DX(nn0939), .F0(\c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_212_) );
      defparam ii0939.CONFIG_DATA = 16'hCACA;
      defparam ii0939.PLACE_LOCATION = "NONE";
      defparam ii0939.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0940 ( .DX(nn0940), .F0(\c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0940.CONFIG_DATA = 16'h35FF;
      defparam ii0940.PLACE_LOCATION = "NONE";
      defparam ii0940.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0941 ( .DX(\a_diny[1]_cal1_u139_mac ), .F0(nn0803), .F1(nn0939), .F2(nn0940), .F3(dummy_abc_213_) );
      defparam ii0941.CONFIG_DATA = 16'h8F8F;
      defparam ii0941.PLACE_LOCATION = "NONE";
      defparam ii0941.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0942 ( .DX(nn0942), .F0(\c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_214_) );
      defparam ii0942.CONFIG_DATA = 16'hCACA;
      defparam ii0942.PLACE_LOCATION = "NONE";
      defparam ii0942.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0943 ( .DX(nn0943), .F0(\c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0943.CONFIG_DATA = 16'h35FF;
      defparam ii0943.PLACE_LOCATION = "NONE";
      defparam ii0943.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0944 ( .DX(\a_diny[1]_cal1_u140_mac ), .F0(nn0803), .F1(nn0942), .F2(nn0943), .F3(dummy_abc_215_) );
      defparam ii0944.CONFIG_DATA = 16'h8F8F;
      defparam ii0944.PLACE_LOCATION = "NONE";
      defparam ii0944.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0945 ( .DX(nn0945), .F0(dummy_123_), .F1(nn0806), .F2(dummy_abc_216_), .F3(dummy_abc_217_) );
      defparam ii0945.CONFIG_DATA = 16'h4444;
      defparam ii0945.PLACE_LOCATION = "NONE";
      defparam ii0945.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0946 ( .DX(nn0946), .F0(\c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0893), .F3(nn0891) );
      defparam ii0946.CONFIG_DATA = 16'h153F;
      defparam ii0946.PLACE_LOCATION = "NONE";
      defparam ii0946.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0947 ( .DX(nn0947), .F0(\c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0946) );
      defparam ii0947.CONFIG_DATA = 16'hDF00;
      defparam ii0947.PLACE_LOCATION = "NONE";
      defparam ii0947.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0948 ( .DX(\a_diny[1]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u139_mac ), .F2(nn0947), .F3(dummy_abc_218_) );
      defparam ii0948.CONFIG_DATA = 16'h8F8F;
      defparam ii0948.PLACE_LOCATION = "NONE";
      defparam ii0948.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0949 ( .DX(nn0949), .F0(\c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0897), .F3(nn0899) );
      defparam ii0949.CONFIG_DATA = 16'h153F;
      defparam ii0949.PLACE_LOCATION = "NONE";
      defparam ii0949.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0950 ( .DX(nn0950), .F0(\c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0898), .F2(nn0949), .F3(dummy_abc_219_) );
      defparam ii0950.CONFIG_DATA = 16'h7070;
      defparam ii0950.PLACE_LOCATION = "NONE";
      defparam ii0950.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0951 ( .DX(\a_diny[1]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u140_mac ), .F2(nn0950), .F3(dummy_abc_220_) );
      defparam ii0951.CONFIG_DATA = 16'h8F8F;
      defparam ii0951.PLACE_LOCATION = "NONE";
      defparam ii0951.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0952 ( .DX(nn0952), .F0(\c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_221_) );
      defparam ii0952.CONFIG_DATA = 16'hCACA;
      defparam ii0952.PLACE_LOCATION = "NONE";
      defparam ii0952.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0953 ( .DX(nn0953), .F0(\c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0953.CONFIG_DATA = 16'h35FF;
      defparam ii0953.PLACE_LOCATION = "NONE";
      defparam ii0953.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0954 ( .DX(\a_diny[1]_cal1_u143_mac ), .F0(nn0803), .F1(nn0952), .F2(nn0953), .F3(dummy_abc_222_) );
      defparam ii0954.CONFIG_DATA = 16'h8F8F;
      defparam ii0954.PLACE_LOCATION = "NONE";
      defparam ii0954.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0955 ( .DX(nn0955), .F0(\c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_223_) );
      defparam ii0955.CONFIG_DATA = 16'hCACA;
      defparam ii0955.PLACE_LOCATION = "NONE";
      defparam ii0955.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0956 ( .DX(nn0956), .F0(\c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0956.CONFIG_DATA = 16'h35FF;
      defparam ii0956.PLACE_LOCATION = "NONE";
      defparam ii0956.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0957 ( .DX(\a_diny[1]_cal1_u144_mac ), .F0(nn0803), .F1(nn0955), .F2(nn0956), .F3(dummy_abc_224_) );
      defparam ii0957.CONFIG_DATA = 16'h8F8F;
      defparam ii0957.PLACE_LOCATION = "NONE";
      defparam ii0957.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0958 ( .DX(nn0958), .F0(\c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0893), .F3(nn0891) );
      defparam ii0958.CONFIG_DATA = 16'h153F;
      defparam ii0958.PLACE_LOCATION = "NONE";
      defparam ii0958.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0959 ( .DX(nn0959), .F0(\c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0958) );
      defparam ii0959.CONFIG_DATA = 16'hDF00;
      defparam ii0959.PLACE_LOCATION = "NONE";
      defparam ii0959.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0960 ( .DX(\a_diny[1]_cal1_u145_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u143_mac ), .F2(nn0959), .F3(dummy_abc_225_) );
      defparam ii0960.CONFIG_DATA = 16'h8F8F;
      defparam ii0960.PLACE_LOCATION = "NONE";
      defparam ii0960.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0961 ( .DX(nn0961), .F0(\c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0897) );
      defparam ii0961.CONFIG_DATA = 16'h135F;
      defparam ii0961.PLACE_LOCATION = "NONE";
      defparam ii0961.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0962 ( .DX(nn0962), .F0(\c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0961) );
      defparam ii0962.CONFIG_DATA = 16'hDF00;
      defparam ii0962.PLACE_LOCATION = "NONE";
      defparam ii0962.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0963 ( .DX(\a_diny[1]_cal1_u146_mac ), .F0(dummy_123_), .F1(\a_diny[1]_cal1_u144_mac ), .F2(nn0962), .F3(dummy_abc_226_) );
      defparam ii0963.CONFIG_DATA = 16'h8F8F;
      defparam ii0963.PLACE_LOCATION = "NONE";
      defparam ii0963.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0964 ( .DX(nn0964), .F0(\c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_227_) );
      defparam ii0964.CONFIG_DATA = 16'hCACA;
      defparam ii0964.PLACE_LOCATION = "NONE";
      defparam ii0964.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0965 ( .DX(nn0965), .F0(\c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0965.CONFIG_DATA = 16'h35FF;
      defparam ii0965.PLACE_LOCATION = "NONE";
      defparam ii0965.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0966 ( .DX(\a_diny[2]_cal1_u135_mac ), .F0(nn0803), .F1(nn0964), .F2(nn0965), .F3(dummy_abc_228_) );
      defparam ii0966.CONFIG_DATA = 16'h8F8F;
      defparam ii0966.PLACE_LOCATION = "NONE";
      defparam ii0966.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0967 ( .DX(nn0967), .F0(\c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_229_) );
      defparam ii0967.CONFIG_DATA = 16'hCACA;
      defparam ii0967.PLACE_LOCATION = "NONE";
      defparam ii0967.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0968 ( .DX(nn0968), .F0(\c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0968.CONFIG_DATA = 16'h35FF;
      defparam ii0968.PLACE_LOCATION = "NONE";
      defparam ii0968.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0969 ( .DX(\a_diny[2]_cal1_u136_mac ), .F0(nn0803), .F1(nn0967), .F2(nn0968), .F3(dummy_abc_230_) );
      defparam ii0969.CONFIG_DATA = 16'h8F8F;
      defparam ii0969.PLACE_LOCATION = "NONE";
      defparam ii0969.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0970 ( .DX(nn0970), .F0(\c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0893) );
      defparam ii0970.CONFIG_DATA = 16'h135F;
      defparam ii0970.PLACE_LOCATION = "NONE";
      defparam ii0970.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0971 ( .DX(nn0971), .F0(\c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0891), .F2(nn0970), .F3(dummy_abc_231_) );
      defparam ii0971.CONFIG_DATA = 16'h7070;
      defparam ii0971.PLACE_LOCATION = "NONE";
      defparam ii0971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0972 ( .DX(\a_diny[2]_cal1_u137_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u135_mac ), .F2(nn0971), .F3(dummy_abc_232_) );
      defparam ii0972.CONFIG_DATA = 16'h8F8F;
      defparam ii0972.PLACE_LOCATION = "NONE";
      defparam ii0972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0973 ( .DX(nn0973), .F0(\c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0897) );
      defparam ii0973.CONFIG_DATA = 16'h135F;
      defparam ii0973.PLACE_LOCATION = "NONE";
      defparam ii0973.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0974 ( .DX(nn0974), .F0(\c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0973) );
      defparam ii0974.CONFIG_DATA = 16'hDF00;
      defparam ii0974.PLACE_LOCATION = "NONE";
      defparam ii0974.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0975 ( .DX(\a_diny[2]_cal1_u138_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u136_mac ), .F2(nn0974), .F3(dummy_abc_233_) );
      defparam ii0975.CONFIG_DATA = 16'h8F8F;
      defparam ii0975.PLACE_LOCATION = "NONE";
      defparam ii0975.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0976 ( .DX(nn0976), .F0(\c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_234_) );
      defparam ii0976.CONFIG_DATA = 16'hCACA;
      defparam ii0976.PLACE_LOCATION = "NONE";
      defparam ii0976.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0977 ( .DX(nn0977), .F0(\c1r2_q[1]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[1]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0977.CONFIG_DATA = 16'h35FF;
      defparam ii0977.PLACE_LOCATION = "NONE";
      defparam ii0977.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0978 ( .DX(\a_diny[2]_cal1_u139_mac ), .F0(nn0803), .F1(nn0976), .F2(nn0977), .F3(dummy_abc_235_) );
      defparam ii0978.CONFIG_DATA = 16'h8F8F;
      defparam ii0978.PLACE_LOCATION = "NONE";
      defparam ii0978.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0979 ( .DX(nn0979), .F0(\c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_236_) );
      defparam ii0979.CONFIG_DATA = 16'h3535;
      defparam ii0979.PLACE_LOCATION = "NONE";
      defparam ii0979.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0980 ( .DX(nn0980), .F0(\c1r2_q[10]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[10]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0980.CONFIG_DATA = 16'h35FF;
      defparam ii0980.PLACE_LOCATION = "NONE";
      defparam ii0980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0981 ( .DX(\a_diny[2]_cal1_u140_mac ), .F0(nn0803), .F1(nn0979), .F2(nn0980), .F3(dummy_abc_237_) );
      defparam ii0981.CONFIG_DATA = 16'h2F2F;
      defparam ii0981.PLACE_LOCATION = "NONE";
      defparam ii0981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0982 ( .DX(nn0982), .F0(\c1r2_q[1]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(\c1r4_q[1]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0893), .F3(nn0891) );
      defparam ii0982.CONFIG_DATA = 16'h153F;
      defparam ii0982.PLACE_LOCATION = "NONE";
      defparam ii0982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0983 ( .DX(nn0983), .F0(\c1r2_q[1]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0982) );
      defparam ii0983.CONFIG_DATA = 16'hDF00;
      defparam ii0983.PLACE_LOCATION = "NONE";
      defparam ii0983.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0984 ( .DX(\a_diny[2]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u139_mac ), .F2(nn0983), .F3(dummy_abc_238_) );
      defparam ii0984.CONFIG_DATA = 16'h8F8F;
      defparam ii0984.PLACE_LOCATION = "NONE";
      defparam ii0984.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0985 ( .DX(nn0985), .F0(\c1r2_q[10]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r2_q[10]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0898), .F3(nn0899) );
      defparam ii0985.CONFIG_DATA = 16'h153F;
      defparam ii0985.PLACE_LOCATION = "NONE";
      defparam ii0985.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0986 ( .DX(nn0986), .F0(\c1r4_q[10]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0897), .F2(nn0985), .F3(dummy_abc_239_) );
      defparam ii0986.CONFIG_DATA = 16'h7070;
      defparam ii0986.PLACE_LOCATION = "NONE";
      defparam ii0986.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0987 ( .DX(\a_diny[2]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u140_mac ), .F2(nn0986), .F3(dummy_abc_240_) );
      defparam ii0987.CONFIG_DATA = 16'h8F8F;
      defparam ii0987.PLACE_LOCATION = "NONE";
      defparam ii0987.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0988 ( .DX(nn0988), .F0(\c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_241_) );
      defparam ii0988.CONFIG_DATA = 16'hCACA;
      defparam ii0988.PLACE_LOCATION = "NONE";
      defparam ii0988.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0989 ( .DX(nn0989), .F0(\c1r1_q[0]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0989.CONFIG_DATA = 16'h35FF;
      defparam ii0989.PLACE_LOCATION = "NONE";
      defparam ii0989.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0990 ( .DX(\a_diny[2]_cal1_u143_mac ), .F0(nn0803), .F1(nn0988), .F2(nn0989), .F3(dummy_abc_242_) );
      defparam ii0990.CONFIG_DATA = 16'h8F8F;
      defparam ii0990.PLACE_LOCATION = "NONE";
      defparam ii0990.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0991 ( .DX(nn0991), .F0(\c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_243_) );
      defparam ii0991.CONFIG_DATA = 16'hCACA;
      defparam ii0991.PLACE_LOCATION = "NONE";
      defparam ii0991.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0992 ( .DX(nn0992), .F0(\c1r1_q[9]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii0992.CONFIG_DATA = 16'h35FF;
      defparam ii0992.PLACE_LOCATION = "NONE";
      defparam ii0992.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0993 ( .DX(\a_diny[2]_cal1_u144_mac ), .F0(nn0803), .F1(nn0991), .F2(nn0992), .F3(dummy_abc_244_) );
      defparam ii0993.CONFIG_DATA = 16'h8F8F;
      defparam ii0993.PLACE_LOCATION = "NONE";
      defparam ii0993.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0994 ( .DX(nn0994), .F0(\c1r1_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0892), .F3(nn0893) );
      defparam ii0994.CONFIG_DATA = 16'h135F;
      defparam ii0994.PLACE_LOCATION = "NONE";
      defparam ii0994.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0995 ( .DX(nn0995), .F0(\c1r1_q[0]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0891), .F2(nn0994), .F3(dummy_abc_245_) );
      defparam ii0995.CONFIG_DATA = 16'h7070;
      defparam ii0995.PLACE_LOCATION = "NONE";
      defparam ii0995.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0996 ( .DX(\a_diny[2]_cal1_u145_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u143_mac ), .F2(nn0995), .F3(dummy_abc_246_) );
      defparam ii0996.CONFIG_DATA = 16'h8F8F;
      defparam ii0996.PLACE_LOCATION = "NONE";
      defparam ii0996.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0997 ( .DX(nn0997), .F0(\c1r1_q[9]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0898), .F3(nn0897) );
      defparam ii0997.CONFIG_DATA = 16'h135F;
      defparam ii0997.PLACE_LOCATION = "NONE";
      defparam ii0997.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0998 ( .DX(nn0998), .F0(\c1r1_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn0997) );
      defparam ii0998.CONFIG_DATA = 16'hDF00;
      defparam ii0998.PLACE_LOCATION = "NONE";
      defparam ii0998.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0999 ( .DX(\a_diny[2]_cal1_u146_mac ), .F0(dummy_123_), .F1(\a_diny[2]_cal1_u144_mac ), .F2(nn0998), .F3(dummy_abc_247_) );
      defparam ii0999.CONFIG_DATA = 16'h8F8F;
      defparam ii0999.PLACE_LOCATION = "NONE";
      defparam ii0999.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1000 ( .DX(nn1000), .F0(\c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_248_) );
      defparam ii1000.CONFIG_DATA = 16'h3535;
      defparam ii1000.PLACE_LOCATION = "NONE";
      defparam ii1000.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1001 ( .DX(nn1001), .F0(\c1r1_q[3]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1001.CONFIG_DATA = 16'h35FF;
      defparam ii1001.PLACE_LOCATION = "NONE";
      defparam ii1001.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1002 ( .DX(\a_diny[3]_cal1_u135_mac ), .F0(nn0803), .F1(nn1000), .F2(nn1001), .F3(dummy_abc_249_) );
      defparam ii1002.CONFIG_DATA = 16'h2F2F;
      defparam ii1002.PLACE_LOCATION = "NONE";
      defparam ii1002.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1003 ( .DX(nn1003), .F0(\c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_250_) );
      defparam ii1003.CONFIG_DATA = 16'h3535;
      defparam ii1003.PLACE_LOCATION = "NONE";
      defparam ii1003.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1004 ( .DX(nn1004), .F0(\c1r1_q[12]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1004.CONFIG_DATA = 16'h35FF;
      defparam ii1004.PLACE_LOCATION = "NONE";
      defparam ii1004.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1005 ( .DX(\a_diny[3]_cal1_u136_mac ), .F0(nn0803), .F1(nn1003), .F2(nn1004), .F3(dummy_abc_251_) );
      defparam ii1005.CONFIG_DATA = 16'h2F2F;
      defparam ii1005.PLACE_LOCATION = "NONE";
      defparam ii1005.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1006 ( .DX(nn1006), .F0(\c1r1_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r1_q[3]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0892), .F3(nn0891) );
      defparam ii1006.CONFIG_DATA = 16'h135F;
      defparam ii1006.PLACE_LOCATION = "NONE";
      defparam ii1006.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1007 ( .DX(nn1007), .F0(\c1r3_q[3]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0893), .F2(nn1006), .F3(dummy_abc_252_) );
      defparam ii1007.CONFIG_DATA = 16'h7070;
      defparam ii1007.PLACE_LOCATION = "NONE";
      defparam ii1007.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1008 ( .DX(\a_diny[3]_cal1_u137_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u135_mac ), .F2(nn1007), .F3(dummy_abc_253_) );
      defparam ii1008.CONFIG_DATA = 16'h8F8F;
      defparam ii1008.PLACE_LOCATION = "NONE";
      defparam ii1008.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1009 ( .DX(nn1009), .F0(\c1r1_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1009.CONFIG_DATA = 16'h153F;
      defparam ii1009.PLACE_LOCATION = "NONE";
      defparam ii1009.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1010 ( .DX(nn1010), .F0(\c1r1_q[12]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0898), .F2(nn1009), .F3(dummy_abc_254_) );
      defparam ii1010.CONFIG_DATA = 16'h7070;
      defparam ii1010.PLACE_LOCATION = "NONE";
      defparam ii1010.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1011 ( .DX(\a_diny[3]_cal1_u138_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u136_mac ), .F2(nn1010), .F3(dummy_abc_255_) );
      defparam ii1011.CONFIG_DATA = 16'h8F8F;
      defparam ii1011.PLACE_LOCATION = "NONE";
      defparam ii1011.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1012 ( .DX(nn1012), .F0(\c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_256_) );
      defparam ii1012.CONFIG_DATA = 16'hCACA;
      defparam ii1012.PLACE_LOCATION = "NONE";
      defparam ii1012.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1013 ( .DX(nn1013), .F0(\c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1013.CONFIG_DATA = 16'h35FF;
      defparam ii1013.PLACE_LOCATION = "NONE";
      defparam ii1013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1014 ( .DX(\a_diny[3]_cal1_u139_mac ), .F0(nn0803), .F1(nn1012), .F2(nn1013), .F3(dummy_abc_257_) );
      defparam ii1014.CONFIG_DATA = 16'h8F8F;
      defparam ii1014.PLACE_LOCATION = "NONE";
      defparam ii1014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1015 ( .DX(nn1015), .F0(\c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_258_) );
      defparam ii1015.CONFIG_DATA = 16'h3535;
      defparam ii1015.PLACE_LOCATION = "NONE";
      defparam ii1015.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1016 ( .DX(nn1016), .F0(\c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1016.CONFIG_DATA = 16'h35FF;
      defparam ii1016.PLACE_LOCATION = "NONE";
      defparam ii1016.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1017 ( .DX(\a_diny[3]_cal1_u140_mac ), .F0(nn0803), .F1(nn1015), .F2(nn1016), .F3(dummy_abc_259_) );
      defparam ii1017.CONFIG_DATA = 16'h2F2F;
      defparam ii1017.PLACE_LOCATION = "NONE";
      defparam ii1017.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1018 ( .DX(nn1018), .F0(\c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0893) );
      defparam ii1018.CONFIG_DATA = 16'h135F;
      defparam ii1018.PLACE_LOCATION = "NONE";
      defparam ii1018.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1019 ( .DX(nn1019), .F0(\c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0891), .F2(nn1018), .F3(dummy_abc_260_) );
      defparam ii1019.CONFIG_DATA = 16'h7070;
      defparam ii1019.PLACE_LOCATION = "NONE";
      defparam ii1019.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1020 ( .DX(\a_diny[3]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u139_mac ), .F2(nn1019), .F3(dummy_abc_261_) );
      defparam ii1020.CONFIG_DATA = 16'h8F8F;
      defparam ii1020.PLACE_LOCATION = "NONE";
      defparam ii1020.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1021 ( .DX(nn1021), .F0(\c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1021.CONFIG_DATA = 16'h153F;
      defparam ii1021.PLACE_LOCATION = "NONE";
      defparam ii1021.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1022 ( .DX(nn1022), .F0(\c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0898), .F2(nn1021), .F3(dummy_abc_262_) );
      defparam ii1022.CONFIG_DATA = 16'h7070;
      defparam ii1022.PLACE_LOCATION = "NONE";
      defparam ii1022.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1023 ( .DX(\a_diny[3]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u140_mac ), .F2(nn1022), .F3(dummy_abc_263_) );
      defparam ii1023.CONFIG_DATA = 16'h8F8F;
      defparam ii1023.PLACE_LOCATION = "NONE";
      defparam ii1023.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1024 ( .DX(nn1024), .F0(\c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_264_) );
      defparam ii1024.CONFIG_DATA = 16'hCACA;
      defparam ii1024.PLACE_LOCATION = "NONE";
      defparam ii1024.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1025 ( .DX(nn1025), .F0(\c1r2_q[0]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[0]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1025.CONFIG_DATA = 16'h35FF;
      defparam ii1025.PLACE_LOCATION = "NONE";
      defparam ii1025.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1026 ( .DX(\a_diny[3]_cal1_u143_mac ), .F0(nn0803), .F1(nn1024), .F2(nn1025), .F3(dummy_abc_265_) );
      defparam ii1026.CONFIG_DATA = 16'h8F8F;
      defparam ii1026.PLACE_LOCATION = "NONE";
      defparam ii1026.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1027 ( .DX(nn1027), .F0(\c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_266_) );
      defparam ii1027.CONFIG_DATA = 16'h3535;
      defparam ii1027.PLACE_LOCATION = "NONE";
      defparam ii1027.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1028 ( .DX(nn1028), .F0(\c1r2_q[9]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[9]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1028.CONFIG_DATA = 16'h35FF;
      defparam ii1028.PLACE_LOCATION = "NONE";
      defparam ii1028.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1029 ( .DX(\a_diny[3]_cal1_u144_mac ), .F0(nn0803), .F1(nn1027), .F2(nn1028), .F3(dummy_abc_267_) );
      defparam ii1029.CONFIG_DATA = 16'h2F2F;
      defparam ii1029.PLACE_LOCATION = "NONE";
      defparam ii1029.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1030 ( .DX(nn1030), .F0(\c1r2_q[0]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(\c1r4_q[0]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0893), .F3(nn0891) );
      defparam ii1030.CONFIG_DATA = 16'h153F;
      defparam ii1030.PLACE_LOCATION = "NONE";
      defparam ii1030.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1031 ( .DX(nn1031), .F0(\c1r2_q[0]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn1030) );
      defparam ii1031.CONFIG_DATA = 16'hDF00;
      defparam ii1031.PLACE_LOCATION = "NONE";
      defparam ii1031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1032 ( .DX(\a_diny[3]_cal1_u145_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u143_mac ), .F2(nn1031), .F3(dummy_abc_268_) );
      defparam ii1032.CONFIG_DATA = 16'h8F8F;
      defparam ii1032.PLACE_LOCATION = "NONE";
      defparam ii1032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1033 ( .DX(nn1033), .F0(\c1r2_q[9]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[9]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1033.CONFIG_DATA = 16'h153F;
      defparam ii1033.PLACE_LOCATION = "NONE";
      defparam ii1033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1034 ( .DX(nn1034), .F0(\c1r2_q[9]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0898), .F2(nn1033), .F3(dummy_abc_269_) );
      defparam ii1034.CONFIG_DATA = 16'h7070;
      defparam ii1034.PLACE_LOCATION = "NONE";
      defparam ii1034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1035 ( .DX(\a_diny[3]_cal1_u146_mac ), .F0(dummy_123_), .F1(\a_diny[3]_cal1_u144_mac ), .F2(nn1034), .F3(dummy_abc_270_) );
      defparam ii1035.CONFIG_DATA = 16'h8F8F;
      defparam ii1035.PLACE_LOCATION = "NONE";
      defparam ii1035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1036 ( .DX(nn1036), .F0(\c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_271_) );
      defparam ii1036.CONFIG_DATA = 16'h3535;
      defparam ii1036.PLACE_LOCATION = "NONE";
      defparam ii1036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1037 ( .DX(nn1037), .F0(\c1r2_q[3]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[3]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1037.CONFIG_DATA = 16'h35FF;
      defparam ii1037.PLACE_LOCATION = "NONE";
      defparam ii1037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1038 ( .DX(\a_diny[4]_cal1_u135_mac ), .F0(nn0803), .F1(nn1036), .F2(nn1037), .F3(dummy_abc_272_) );
      defparam ii1038.CONFIG_DATA = 16'h2F2F;
      defparam ii1038.PLACE_LOCATION = "NONE";
      defparam ii1038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1039 ( .DX(nn1039), .F0(\c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_273_) );
      defparam ii1039.CONFIG_DATA = 16'h3535;
      defparam ii1039.PLACE_LOCATION = "NONE";
      defparam ii1039.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1040 ( .DX(nn1040), .F0(\c1r2_q[12]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r4_q[12]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1040.CONFIG_DATA = 16'h35FF;
      defparam ii1040.PLACE_LOCATION = "NONE";
      defparam ii1040.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1041 ( .DX(\a_diny[4]_cal1_u136_mac ), .F0(nn0803), .F1(nn1039), .F2(nn1040), .F3(dummy_abc_274_) );
      defparam ii1041.CONFIG_DATA = 16'h2F2F;
      defparam ii1041.PLACE_LOCATION = "NONE";
      defparam ii1041.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1042 ( .DX(nn1042), .F0(\c1r2_q[3]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r2_q[3]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0892), .F3(nn0891) );
      defparam ii1042.CONFIG_DATA = 16'h135F;
      defparam ii1042.PLACE_LOCATION = "NONE";
      defparam ii1042.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1043 ( .DX(nn1043), .F0(\c1r4_q[3]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0893), .F2(nn1042), .F3(dummy_abc_275_) );
      defparam ii1043.CONFIG_DATA = 16'h7070;
      defparam ii1043.PLACE_LOCATION = "NONE";
      defparam ii1043.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1044 ( .DX(\a_diny[4]_cal1_u137_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u135_mac ), .F2(nn1043), .F3(dummy_abc_276_) );
      defparam ii1044.CONFIG_DATA = 16'h8F8F;
      defparam ii1044.PLACE_LOCATION = "NONE";
      defparam ii1044.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1045 ( .DX(nn1045), .F0(\c1r2_q[12]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r4_q[12]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1045.CONFIG_DATA = 16'h153F;
      defparam ii1045.PLACE_LOCATION = "NONE";
      defparam ii1045.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1046 ( .DX(nn1046), .F0(\c1r2_q[12]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0898), .F2(nn1045), .F3(dummy_abc_277_) );
      defparam ii1046.CONFIG_DATA = 16'h7070;
      defparam ii1046.PLACE_LOCATION = "NONE";
      defparam ii1046.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1047 ( .DX(\a_diny[4]_cal1_u138_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u136_mac ), .F2(nn1046), .F3(dummy_abc_278_) );
      defparam ii1047.CONFIG_DATA = 16'h8F8F;
      defparam ii1047.PLACE_LOCATION = "NONE";
      defparam ii1047.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1048 ( .DX(nn1048), .F0(\c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_279_) );
      defparam ii1048.CONFIG_DATA = 16'hCACA;
      defparam ii1048.PLACE_LOCATION = "NONE";
      defparam ii1048.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1049 ( .DX(nn1049), .F0(\c1r2_q[2]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1049.CONFIG_DATA = 16'h35FF;
      defparam ii1049.PLACE_LOCATION = "NONE";
      defparam ii1049.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1050 ( .DX(\a_diny[4]_cal1_u139_mac ), .F0(nn0803), .F1(nn1048), .F2(nn1049), .F3(dummy_abc_280_) );
      defparam ii1050.CONFIG_DATA = 16'h8F8F;
      defparam ii1050.PLACE_LOCATION = "NONE";
      defparam ii1050.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1051 ( .DX(nn1051), .F0(\c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_281_) );
      defparam ii1051.CONFIG_DATA = 16'hCACA;
      defparam ii1051.PLACE_LOCATION = "NONE";
      defparam ii1051.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1052 ( .DX(nn1052), .F0(\c1r2_q[11]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1052.CONFIG_DATA = 16'h35FF;
      defparam ii1052.PLACE_LOCATION = "NONE";
      defparam ii1052.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1053 ( .DX(\a_diny[4]_cal1_u140_mac ), .F0(nn0803), .F1(nn1051), .F2(nn1052), .F3(dummy_abc_282_) );
      defparam ii1053.CONFIG_DATA = 16'h8F8F;
      defparam ii1053.PLACE_LOCATION = "NONE";
      defparam ii1053.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1054 ( .DX(nn1054), .F0(\c1r2_q[2]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0893), .F3(nn0891) );
      defparam ii1054.CONFIG_DATA = 16'h153F;
      defparam ii1054.PLACE_LOCATION = "NONE";
      defparam ii1054.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1055 ( .DX(nn1055), .F0(\c1r2_q[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn1054) );
      defparam ii1055.CONFIG_DATA = 16'hDF00;
      defparam ii1055.PLACE_LOCATION = "NONE";
      defparam ii1055.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1056 ( .DX(\a_diny[4]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u139_mac ), .F2(nn1055), .F3(dummy_abc_283_) );
      defparam ii1056.CONFIG_DATA = 16'h8F8F;
      defparam ii1056.PLACE_LOCATION = "NONE";
      defparam ii1056.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1057 ( .DX(nn1057), .F0(\c1r2_q[11]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0898), .F3(nn0897) );
      defparam ii1057.CONFIG_DATA = 16'h135F;
      defparam ii1057.PLACE_LOCATION = "NONE";
      defparam ii1057.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1058 ( .DX(nn1058), .F0(\c1r2_q[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn1057) );
      defparam ii1058.CONFIG_DATA = 16'hDF00;
      defparam ii1058.PLACE_LOCATION = "NONE";
      defparam ii1058.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1059 ( .DX(\a_diny[4]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u140_mac ), .F2(nn1058), .F3(dummy_abc_284_) );
      defparam ii1059.CONFIG_DATA = 16'h8F8F;
      defparam ii1059.PLACE_LOCATION = "NONE";
      defparam ii1059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1060 ( .DX(nn1060), .F0(\c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_285_) );
      defparam ii1060.CONFIG_DATA = 16'hCACA;
      defparam ii1060.PLACE_LOCATION = "NONE";
      defparam ii1060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1061 ( .DX(nn1061), .F0(\c1r1_q[1]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1061.CONFIG_DATA = 16'h35FF;
      defparam ii1061.PLACE_LOCATION = "NONE";
      defparam ii1061.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1062 ( .DX(\a_diny[4]_cal1_u143_mac ), .F0(nn0803), .F1(nn1060), .F2(nn1061), .F3(dummy_abc_286_) );
      defparam ii1062.CONFIG_DATA = 16'h8F8F;
      defparam ii1062.PLACE_LOCATION = "NONE";
      defparam ii1062.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1063 ( .DX(nn1063), .F0(\c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_287_) );
      defparam ii1063.CONFIG_DATA = 16'h3535;
      defparam ii1063.PLACE_LOCATION = "NONE";
      defparam ii1063.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1064 ( .DX(nn1064), .F0(\c1r1_q[10]_fifo1_ram_inst_3_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_3_u_emb18k_0 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1064.CONFIG_DATA = 16'h35FF;
      defparam ii1064.PLACE_LOCATION = "NONE";
      defparam ii1064.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1065 ( .DX(\a_diny[4]_cal1_u144_mac ), .F0(nn0803), .F1(nn1063), .F2(nn1064), .F3(dummy_abc_288_) );
      defparam ii1065.CONFIG_DATA = 16'h2F2F;
      defparam ii1065.PLACE_LOCATION = "NONE";
      defparam ii1065.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1066 ( .DX(nn1066), .F0(\c1r1_q[1]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r1_q[1]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0892), .F3(nn0891) );
      defparam ii1066.CONFIG_DATA = 16'h135F;
      defparam ii1066.PLACE_LOCATION = "NONE";
      defparam ii1066.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1067 ( .DX(nn1067), .F0(\c1r3_q[1]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0893), .F2(nn1066), .F3(dummy_abc_289_) );
      defparam ii1067.CONFIG_DATA = 16'h7070;
      defparam ii1067.PLACE_LOCATION = "NONE";
      defparam ii1067.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1068 ( .DX(\a_diny[4]_cal1_u145_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u143_mac ), .F2(nn1067), .F3(dummy_abc_290_) );
      defparam ii1068.CONFIG_DATA = 16'h8F8F;
      defparam ii1068.PLACE_LOCATION = "NONE";
      defparam ii1068.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1069 ( .DX(nn1069), .F0(\c1r1_q[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1_u_emb18k_0 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1069.CONFIG_DATA = 16'h153F;
      defparam ii1069.PLACE_LOCATION = "NONE";
      defparam ii1069.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1070 ( .DX(nn1070), .F0(\c1r1_q[10]_fifo1_ram_inst_1_u_emb18k_0 ), .F1(nn0898), .F2(nn1069), .F3(dummy_abc_291_) );
      defparam ii1070.CONFIG_DATA = 16'h7070;
      defparam ii1070.PLACE_LOCATION = "NONE";
      defparam ii1070.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1071 ( .DX(\a_diny[4]_cal1_u146_mac ), .F0(dummy_123_), .F1(\a_diny[4]_cal1_u144_mac ), .F2(nn1070), .F3(dummy_abc_292_) );
      defparam ii1071.CONFIG_DATA = 16'h8F8F;
      defparam ii1071.PLACE_LOCATION = "NONE";
      defparam ii1071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1072 ( .DX(nn1072), .F0(\c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_293_) );
      defparam ii1072.CONFIG_DATA = 16'hCACA;
      defparam ii1072.PLACE_LOCATION = "NONE";
      defparam ii1072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1073 ( .DX(nn1073), .F0(\c1r1_q[2]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_aa_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1073.CONFIG_DATA = 16'h35FF;
      defparam ii1073.PLACE_LOCATION = "NONE";
      defparam ii1073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1074 ( .DX(\a_diny[5]_cal1_u139_mac ), .F0(nn0803), .F1(nn1072), .F2(nn1073), .F3(dummy_abc_294_) );
      defparam ii1074.CONFIG_DATA = 16'h8F8F;
      defparam ii1074.PLACE_LOCATION = "NONE";
      defparam ii1074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1075 ( .DX(nn1075), .F0(\c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F2(\fifo1_ram_inst_0_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_295_) );
      defparam ii1075.CONFIG_DATA = 16'h3535;
      defparam ii1075.PLACE_LOCATION = "NONE";
      defparam ii1075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1076 ( .DX(nn1076), .F0(\c1r1_q[11]_fifo1_ram_inst_3_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_3_u_emb18k_1 ), .F2(\fifo1_ram_inst_3_ab_reg__reg[0]|Q_net ), .F3(nn0806) );
      defparam ii1076.CONFIG_DATA = 16'h35FF;
      defparam ii1076.PLACE_LOCATION = "NONE";
      defparam ii1076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1077 ( .DX(\a_diny[5]_cal1_u140_mac ), .F0(nn0803), .F1(nn1075), .F2(nn1076), .F3(dummy_abc_296_) );
      defparam ii1077.CONFIG_DATA = 16'h2F2F;
      defparam ii1077.PLACE_LOCATION = "NONE";
      defparam ii1077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1078 ( .DX(nn1078), .F0(\c1r1_q[2]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0893), .F3(nn0891) );
      defparam ii1078.CONFIG_DATA = 16'h153F;
      defparam ii1078.PLACE_LOCATION = "NONE";
      defparam ii1078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1079 ( .DX(nn1079), .F0(\c1r1_q[2]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\fifo1_ram_inst_0_aa_reg__reg[0]|Q_net ), .F2(nn0945), .F3(nn1078) );
      defparam ii1079.CONFIG_DATA = 16'hDF00;
      defparam ii1079.PLACE_LOCATION = "NONE";
      defparam ii1079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1080 ( .DX(\a_diny[5]_cal1_u141_mac ), .F0(dummy_123_), .F1(\a_diny[5]_cal1_u139_mac ), .F2(nn1079), .F3(dummy_abc_297_) );
      defparam ii1080.CONFIG_DATA = 16'h8F8F;
      defparam ii1080.PLACE_LOCATION = "NONE";
      defparam ii1080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1081 ( .DX(nn1081), .F0(\c1r1_q[11]_fifo1_ram_inst_0_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1_u_emb18k_1 ), .F2(nn0897), .F3(nn0899) );
      defparam ii1081.CONFIG_DATA = 16'h153F;
      defparam ii1081.PLACE_LOCATION = "NONE";
      defparam ii1081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1082 ( .DX(nn1082), .F0(\c1r1_q[11]_fifo1_ram_inst_1_u_emb18k_1 ), .F1(nn0898), .F2(nn1081), .F3(dummy_abc_298_) );
      defparam ii1082.CONFIG_DATA = 16'h7070;
      defparam ii1082.PLACE_LOCATION = "NONE";
      defparam ii1082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1083 ( .DX(\a_diny[5]_cal1_u142_mac ), .F0(dummy_123_), .F1(\a_diny[5]_cal1_u140_mac ), .F2(nn1082), .F3(dummy_abc_299_) );
      defparam ii1083.CONFIG_DATA = 16'h8F8F;
      defparam ii1083.PLACE_LOCATION = "NONE";
      defparam ii1083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1084 ( .DX(u6796_O), .F0(rst), .F1(u4510_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(dummy_abc_300_) );
      defparam ii1084.CONFIG_DATA = 16'hEAEA;
      defparam ii1084.PLACE_LOCATION = "NONE";
      defparam ii1084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1085 ( .DX(u6789_Y), .F0(rst), .F1(u6810_IN), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(nn0801) );
      defparam ii1085.CONFIG_DATA = 16'h1441;
      defparam ii1085.PLACE_LOCATION = "NONE";
      defparam ii1085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1086 ( .DX(nn1086), .F0(u6810_D0), .F1(u6810_I0_3_), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(u6789_Y) );
      defparam ii1086.CONFIG_DATA = 16'hC535;
      defparam ii1086.PLACE_LOCATION = "NONE";
      defparam ii1086.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1087 ( .DX(nn1087), .F0(u6810_I0), .F1(u6810_I0_0_), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(u6789_Y) );
      defparam ii1087.CONFIG_DATA = 16'h5553;
      defparam ii1087.PLACE_LOCATION = "NONE";
      defparam ii1087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1088 ( .DX(nn1088), .F0(\cal1_jmp2Normal__reg|Q_net ), .F1(nn0801), .F2(nn1086), .F3(nn1087) );
      defparam ii1088.CONFIG_DATA = 16'hC8FB;
      defparam ii1088.PLACE_LOCATION = "NONE";
      defparam ii1088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1089 ( .DX(nn1089), .F0(rst), .F1(u6810_I0_0_), .F2(nn0801), .F3(dummy_abc_301_) );
      defparam ii1089.CONFIG_DATA = 16'h1010;
      defparam ii1089.PLACE_LOCATION = "NONE";
      defparam ii1089.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1090 ( .DX(nn1090), .F0(u6810_I0), .F1(\inputctrl1_jmp__reg|Q_net ), .F2(u6789_Y), .F3(nn1089) );
      defparam ii1090.CONFIG_DATA = 16'h80BF;
      defparam ii1090.PLACE_LOCATION = "NONE";
      defparam ii1090.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1091 ( .DX(u3634_OUT), .F0(rst), .F1(\cal1_jmp2Normal__reg|Q_net ), .F2(nn1088), .F3(nn1090) );
      defparam ii1091.CONFIG_DATA = 16'hFA32;
      defparam ii1091.PLACE_LOCATION = "NONE";
      defparam ii1091.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1092 ( .DX(nn1092), .F0(nn0802), .F1(u3634_OUT), .F2(u6796_O), .F3(dummy_abc_302_) );
      defparam ii1092.CONFIG_DATA = 16'h0808;
      defparam ii1092.PLACE_LOCATION = "NONE";
      defparam ii1092.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1093 ( .DX(\c1r1_aa[10]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1093.CONFIG_DATA = 16'h00CA;
      defparam ii1093.PLACE_LOCATION = "NONE";
      defparam ii1093.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1094 ( .DX(nn1094), .F0(rst), .F1(u4510_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(dummy_abc_303_) );
      defparam ii1094.CONFIG_DATA = 16'h4040;
      defparam ii1094.PLACE_LOCATION = "NONE";
      defparam ii1094.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1095 ( .DX(nn1095), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1095.CONFIG_DATA = 16'h33F5;
      defparam ii1095.PLACE_LOCATION = "NONE";
      defparam ii1095.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1096 ( .DX(u3662_O), .F0(rst), .F1(nn0805), .F2(dummy_abc_304_), .F3(dummy_abc_305_) );
      defparam ii1096.CONFIG_DATA = 16'h4444;
      defparam ii1096.PLACE_LOCATION = "NONE";
      defparam ii1096.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1097 ( .DX(\c1r1_aa[10]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(nn1094), .F2(nn1095), .F3(u3662_O) );
      defparam ii1097.CONFIG_DATA = 16'h2F0F;
      defparam ii1097.PLACE_LOCATION = "NONE";
      defparam ii1097.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1098 ( .DX(u3672_O), .F0(rst), .F1(\cal1_jmp2Normal__reg|Q_net ), .F2(nn0801), .F3(nn0802) );
      defparam ii1098.CONFIG_DATA = 16'h0045;
      defparam ii1098.PLACE_LOCATION = "NONE";
      defparam ii1098.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1099 ( .DX(\c1r1_aa[10]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(nn1094), .F2(nn1095), .F3(u3672_O) );
      defparam ii1099.CONFIG_DATA = 16'h2F0F;
      defparam ii1099.PLACE_LOCATION = "NONE";
      defparam ii1099.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1100 ( .DX(\c1r1_aa[11]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1100.CONFIG_DATA = 16'h00CA;
      defparam ii1100.PLACE_LOCATION = "NONE";
      defparam ii1100.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1101 ( .DX(nn1101), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1101.CONFIG_DATA = 16'h33F5;
      defparam ii1101.PLACE_LOCATION = "NONE";
      defparam ii1101.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1102 ( .DX(\c1r1_aa[11]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1101) );
      defparam ii1102.CONFIG_DATA = 16'h20FF;
      defparam ii1102.PLACE_LOCATION = "NONE";
      defparam ii1102.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1103 ( .DX(\c1r1_aa[11]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1101) );
      defparam ii1103.CONFIG_DATA = 16'h20FF;
      defparam ii1103.PLACE_LOCATION = "NONE";
      defparam ii1103.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1104 ( .DX(\c1r1_aa[2]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1104.CONFIG_DATA = 16'h00CA;
      defparam ii1104.PLACE_LOCATION = "NONE";
      defparam ii1104.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1105 ( .DX(nn1105), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1105.CONFIG_DATA = 16'h33F5;
      defparam ii1105.PLACE_LOCATION = "NONE";
      defparam ii1105.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1106 ( .DX(\c1r1_aa[2]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1105) );
      defparam ii1106.CONFIG_DATA = 16'h20FF;
      defparam ii1106.PLACE_LOCATION = "NONE";
      defparam ii1106.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1107 ( .DX(\c1r1_aa[2]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1105) );
      defparam ii1107.CONFIG_DATA = 16'h20FF;
      defparam ii1107.PLACE_LOCATION = "NONE";
      defparam ii1107.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1108 ( .DX(\c1r1_aa[3]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1108.CONFIG_DATA = 16'h00CA;
      defparam ii1108.PLACE_LOCATION = "NONE";
      defparam ii1108.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1109 ( .DX(nn1109), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1109.CONFIG_DATA = 16'h33F5;
      defparam ii1109.PLACE_LOCATION = "NONE";
      defparam ii1109.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1110 ( .DX(\c1r1_aa[3]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1109) );
      defparam ii1110.CONFIG_DATA = 16'h20FF;
      defparam ii1110.PLACE_LOCATION = "NONE";
      defparam ii1110.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1111 ( .DX(\c1r1_aa[3]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1109) );
      defparam ii1111.CONFIG_DATA = 16'h20FF;
      defparam ii1111.PLACE_LOCATION = "NONE";
      defparam ii1111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1112 ( .DX(\c1r1_aa[4]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1112.CONFIG_DATA = 16'h00CA;
      defparam ii1112.PLACE_LOCATION = "NONE";
      defparam ii1112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1113 ( .DX(nn1113), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1113.CONFIG_DATA = 16'h33F5;
      defparam ii1113.PLACE_LOCATION = "NONE";
      defparam ii1113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1114 ( .DX(\c1r1_aa[4]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1113) );
      defparam ii1114.CONFIG_DATA = 16'h20FF;
      defparam ii1114.PLACE_LOCATION = "NONE";
      defparam ii1114.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1115 ( .DX(\c1r1_aa[4]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1113) );
      defparam ii1115.CONFIG_DATA = 16'h20FF;
      defparam ii1115.PLACE_LOCATION = "NONE";
      defparam ii1115.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1116 ( .DX(\c1r1_aa[5]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1116.CONFIG_DATA = 16'h00CA;
      defparam ii1116.PLACE_LOCATION = "NONE";
      defparam ii1116.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1117 ( .DX(nn1117), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1117.CONFIG_DATA = 16'h33F5;
      defparam ii1117.PLACE_LOCATION = "NONE";
      defparam ii1117.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1118 ( .DX(\c1r1_aa[5]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1117) );
      defparam ii1118.CONFIG_DATA = 16'h20FF;
      defparam ii1118.PLACE_LOCATION = "NONE";
      defparam ii1118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1119 ( .DX(\c1r1_aa[5]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1117) );
      defparam ii1119.CONFIG_DATA = 16'h20FF;
      defparam ii1119.PLACE_LOCATION = "NONE";
      defparam ii1119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1120 ( .DX(\c1r1_aa[6]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1120.CONFIG_DATA = 16'h00CA;
      defparam ii1120.PLACE_LOCATION = "NONE";
      defparam ii1120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1121 ( .DX(nn1121), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1121.CONFIG_DATA = 16'h33F5;
      defparam ii1121.PLACE_LOCATION = "NONE";
      defparam ii1121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1122 ( .DX(\c1r1_aa[6]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1121) );
      defparam ii1122.CONFIG_DATA = 16'h20FF;
      defparam ii1122.PLACE_LOCATION = "NONE";
      defparam ii1122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1123 ( .DX(\c1r1_aa[6]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1121) );
      defparam ii1123.CONFIG_DATA = 16'h20FF;
      defparam ii1123.PLACE_LOCATION = "NONE";
      defparam ii1123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1124 ( .DX(\c1r1_aa[7]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1124.CONFIG_DATA = 16'h00CA;
      defparam ii1124.PLACE_LOCATION = "NONE";
      defparam ii1124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1125 ( .DX(nn1125), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1125.CONFIG_DATA = 16'h33F5;
      defparam ii1125.PLACE_LOCATION = "NONE";
      defparam ii1125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1126 ( .DX(\c1r1_aa[7]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1125) );
      defparam ii1126.CONFIG_DATA = 16'h20FF;
      defparam ii1126.PLACE_LOCATION = "NONE";
      defparam ii1126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1127 ( .DX(\c1r1_aa[7]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1125) );
      defparam ii1127.CONFIG_DATA = 16'h20FF;
      defparam ii1127.PLACE_LOCATION = "NONE";
      defparam ii1127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1128 ( .DX(\c1r1_aa[8]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1128.CONFIG_DATA = 16'h00CA;
      defparam ii1128.PLACE_LOCATION = "NONE";
      defparam ii1128.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1129 ( .DX(nn1129), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1129.CONFIG_DATA = 16'h33F5;
      defparam ii1129.PLACE_LOCATION = "NONE";
      defparam ii1129.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1130 ( .DX(\c1r1_aa[8]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1129) );
      defparam ii1130.CONFIG_DATA = 16'h20FF;
      defparam ii1130.PLACE_LOCATION = "NONE";
      defparam ii1130.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1131 ( .DX(\c1r1_aa[8]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1129) );
      defparam ii1131.CONFIG_DATA = 16'h20FF;
      defparam ii1131.PLACE_LOCATION = "NONE";
      defparam ii1131.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1132 ( .DX(\c1r1_aa[9]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1132.CONFIG_DATA = 16'h00CA;
      defparam ii1132.PLACE_LOCATION = "NONE";
      defparam ii1132.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1133 ( .DX(nn1133), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1133.CONFIG_DATA = 16'h33F5;
      defparam ii1133.PLACE_LOCATION = "NONE";
      defparam ii1133.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1134 ( .DX(\c1r1_aa[9]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1133) );
      defparam ii1134.CONFIG_DATA = 16'h20FF;
      defparam ii1134.PLACE_LOCATION = "NONE";
      defparam ii1134.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1135 ( .DX(\c1r1_aa[9]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1133) );
      defparam ii1135.CONFIG_DATA = 16'h20FF;
      defparam ii1135.PLACE_LOCATION = "NONE";
      defparam ii1135.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1136 ( .DX(nn1136), .F0(\cal1_u__reg[6]|Q_net ), .F1(nn0812), .F2(dummy_abc_306_), .F3(dummy_abc_307_) );
      defparam ii1136.CONFIG_DATA = 16'h6666;
      defparam ii1136.PLACE_LOCATION = "NONE";
      defparam ii1136.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1137 ( .DX(nn1137), .F0(\cal1_u__reg[7]|Q_net ), .F1(\u3_XORCI_1|SUM_net ), .F2(dummy_abc_308_), .F3(dummy_abc_309_) );
      defparam ii1137.CONFIG_DATA = 16'h9999;
      defparam ii1137.PLACE_LOCATION = "NONE";
      defparam ii1137.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1138 ( .DX(nn1138), .F0(\cal1_u__reg[8]|Q_net ), .F1(\u3_XORCI_2|SUM_net ), .F2(dummy_abc_310_), .F3(dummy_abc_311_) );
      defparam ii1138.CONFIG_DATA = 16'h9999;
      defparam ii1138.PLACE_LOCATION = "NONE";
      defparam ii1138.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1139 ( .DX(nn1139), .F0(\cal1_u__reg[9]|Q_net ), .F1(\u3_XORCI_3|SUM_net ), .F2(dummy_abc_312_), .F3(dummy_abc_313_) );
      defparam ii1139.CONFIG_DATA = 16'h9999;
      defparam ii1139.PLACE_LOCATION = "NONE";
      defparam ii1139.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1140 ( .DX(nn1140), .F0(\cal1_u__reg[10]|Q_net ), .F1(\u3_XORCI_4|SUM_net ), .F2(dummy_abc_314_), .F3(dummy_abc_315_) );
      defparam ii1140.CONFIG_DATA = 16'h9999;
      defparam ii1140.PLACE_LOCATION = "NONE";
      defparam ii1140.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1141 ( .DX(nn1141), .F0(\cal1_u__reg[11]|Q_net ), .F1(\u3_XORCI_5|SUM_net ), .F2(dummy_abc_316_), .F3(dummy_abc_317_) );
      defparam ii1141.CONFIG_DATA = 16'h9999;
      defparam ii1141.PLACE_LOCATION = "NONE";
      defparam ii1141.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1142 ( .DX(nn1142), .F0(\cal1_u__reg[12]|Q_net ), .F1(\u3_XORCI_6|SUM_net ), .F2(dummy_abc_318_), .F3(dummy_abc_319_) );
      defparam ii1142.CONFIG_DATA = 16'h9999;
      defparam ii1142.PLACE_LOCATION = "NONE";
      defparam ii1142.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1143 ( .DX(nn1143), .F0(\cal1_u__reg[13]|Q_net ), .F1(\u3_XORCI_7|SUM_net ), .F2(dummy_abc_320_), .F3(dummy_abc_321_) );
      defparam ii1143.CONFIG_DATA = 16'h9999;
      defparam ii1143.PLACE_LOCATION = "NONE";
      defparam ii1143.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1144 ( .DX(nn1144), .F0(\cal1_u__reg[14]|Q_net ), .F1(\u3_XORCI_8|SUM_net ), .F2(dummy_abc_322_), .F3(dummy_abc_323_) );
      defparam ii1144.CONFIG_DATA = 16'h9999;
      defparam ii1144.PLACE_LOCATION = "NONE";
      defparam ii1144.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1145 ( .DX(nn1145), .F0(\cal1_u__reg[15]|Q_net ), .F1(\u3_XORCI_9|SUM_net ), .F2(dummy_abc_324_), .F3(dummy_abc_325_) );
      defparam ii1145.CONFIG_DATA = 16'h9999;
      defparam ii1145.PLACE_LOCATION = "NONE";
      defparam ii1145.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1146 ( .DX(nn1146), .F0(\cal1_u__reg[16]|Q_net ), .F1(\u3_XORCI_10|SUM_net ), .F2(dummy_abc_326_), .F3(dummy_abc_327_) );
      defparam ii1146.CONFIG_DATA = 16'h9999;
      defparam ii1146.PLACE_LOCATION = "NONE";
      defparam ii1146.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1147 ( .DX(nn1147), .F0(dummy_abc_328_), .F1(dummy_abc_329_), .F2(dummy_abc_330_), .F3(dummy_abc_331_) );
      defparam ii1147.CONFIG_DATA = 16'hFFFF;
      defparam ii1147.PLACE_LOCATION = "NONE";
      defparam ii1147.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_7_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \cal1_u__reg[16]|Q_net , 
              \cal1_u__reg[15]|Q_net , \cal1_u__reg[14]|Q_net , \cal1_u__reg[13]|Q_net , 
              \cal1_u__reg[12]|Q_net , \cal1_u__reg[11]|Q_net , \cal1_u__reg[10]|Q_net , 
              \cal1_u__reg[9]|Q_net , \cal1_u__reg[8]|Q_net , \cal1_u__reg[7]|Q_net , 
              \cal1_u__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_52_ ), 
        .DX( {nn1147, nn1146, nn1145, nn1144, nn1143, nn1142, nn1141, nn1140, 
              nn1139, nn1138, nn1137, nn1136} ), 
        .SUM( {\cal1_u61_XORCI_11|SUM_net , dummy_53_, dummy_54_, dummy_55_, 
              dummy_56_, dummy_57_, dummy_58_, dummy_59_, dummy_60_, dummy_61_, 
              dummy_62_, dummy_63_} )
      );
    CS_LUT4_PRIM ii1162 ( .DX(nn1162), .F0(dummy_52_), .F1(dummy_abc_332_), .F2(dummy_abc_333_), .F3(dummy_abc_334_) );
      defparam ii1162.CONFIG_DATA = 16'h5555;
      defparam ii1162.PLACE_LOCATION = "NONE";
      defparam ii1162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1163 ( .DX(nn1163), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(dummy_52_), .F2(dummy_abc_335_), .F3(dummy_abc_336_) );
      defparam ii1163.CONFIG_DATA = 16'h9999;
      defparam ii1163.PLACE_LOCATION = "NONE";
      defparam ii1163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1164 ( .DX(nn1164), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(dummy_abc_337_), .F2(dummy_abc_338_), .F3(dummy_abc_339_) );
      defparam ii1164.CONFIG_DATA = 16'hAAAA;
      defparam ii1164.PLACE_LOCATION = "NONE";
      defparam ii1164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1165 ( .DX(nn1165), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(dummy_abc_340_), .F2(dummy_abc_341_), .F3(dummy_abc_342_) );
      defparam ii1165.CONFIG_DATA = 16'hAAAA;
      defparam ii1165.PLACE_LOCATION = "NONE";
      defparam ii1165.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1166 ( .DX(nn1166), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(dummy_abc_343_), .F2(dummy_abc_344_), .F3(dummy_abc_345_) );
      defparam ii1166.CONFIG_DATA = 16'hAAAA;
      defparam ii1166.PLACE_LOCATION = "NONE";
      defparam ii1166.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1167 ( .DX(nn1167), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(dummy_abc_346_), .F2(dummy_abc_347_), .F3(dummy_abc_348_) );
      defparam ii1167.CONFIG_DATA = 16'hAAAA;
      defparam ii1167.PLACE_LOCATION = "NONE";
      defparam ii1167.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1168 ( .DX(nn1168), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(dummy_abc_349_), .F2(dummy_abc_350_), .F3(dummy_abc_351_) );
      defparam ii1168.CONFIG_DATA = 16'hAAAA;
      defparam ii1168.PLACE_LOCATION = "NONE";
      defparam ii1168.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1169 ( .DX(nn1169), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(dummy_abc_352_), .F2(dummy_abc_353_), .F3(dummy_abc_354_) );
      defparam ii1169.CONFIG_DATA = 16'hAAAA;
      defparam ii1169.PLACE_LOCATION = "NONE";
      defparam ii1169.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1170 ( .DX(nn1170), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(dummy_abc_355_), .F2(dummy_abc_356_), .F3(dummy_abc_357_) );
      defparam ii1170.CONFIG_DATA = 16'hAAAA;
      defparam ii1170.PLACE_LOCATION = "NONE";
      defparam ii1170.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1171 ( .DX(nn1171), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(dummy_abc_358_), .F2(dummy_abc_359_), .F3(dummy_abc_360_) );
      defparam ii1171.CONFIG_DATA = 16'hAAAA;
      defparam ii1171.PLACE_LOCATION = "NONE";
      defparam ii1171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1172 ( .DX(nn1172), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(dummy_abc_361_), .F2(dummy_abc_362_), .F3(dummy_abc_363_) );
      defparam ii1172.CONFIG_DATA = 16'hAAAA;
      defparam ii1172.PLACE_LOCATION = "NONE";
      defparam ii1172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1173 ( .DX(nn1173), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(dummy_abc_364_), .F2(dummy_abc_365_), .F3(dummy_abc_366_) );
      defparam ii1173.CONFIG_DATA = 16'hAAAA;
      defparam ii1173.PLACE_LOCATION = "NONE";
      defparam ii1173.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11 ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1162} ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_12_ ), 
        .DX( {nn1173, nn1172, nn1171, nn1170, nn1169, nn1168, nn1167, nn1166, 
              nn1165, nn1164, nn1163} ), 
        .SUM( {\cal1_u129_XORCI_10|SUM_net , \cal1_u129_XORCI_9|SUM_net , 
              \cal1_u129_XORCI_8|SUM_net , \cal1_u129_XORCI_7|SUM_net , \cal1_u129_XORCI_6|SUM_net , 
              \cal1_u129_XORCI_5|SUM_net , \cal1_u129_XORCI_4|SUM_net , \cal1_u129_XORCI_3|SUM_net , 
              \cal1_u129_XORCI_2|SUM_net , \cal1_u129_XORCI_1|SUM_net , \cal1_u129_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1187 ( .DX(c1r1_clka_fifo1_ram_inst_0_u_emb18k_0), .F0(clka), .F1(clkb), .F2(u6796_O), .F3(dummy_abc_367_) );
      defparam ii1187.CONFIG_DATA = 16'hACAC;
      defparam ii1187.PLACE_LOCATION = "NONE";
      defparam ii1187.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1188 ( .DX(c1r1_clka_fifo1_ram_inst_1_u_emb18k_0), .F0(clka), .F1(clkb), .F2(nn1094), .F3(dummy_abc_368_) );
      defparam ii1188.CONFIG_DATA = 16'hACAC;
      defparam ii1188.PLACE_LOCATION = "NONE";
      defparam ii1188.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1189 ( .DX(dOut[0]), .F0(\a_mac_out[6]_cal1_u143_mac ), .F1(\a_mac_out[6]_cal1_u144_mac ), .F2(\a_mac_out[6]_cal1_u145_mac ), .F3(\a_mac_out[6]_cal1_u146_mac ) );
      defparam ii1189.CONFIG_DATA = 16'h6996;
      defparam ii1189.PLACE_LOCATION = "NONE";
      defparam ii1189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1190 ( .DX(nn1190), .F0(\a_mac_out[6]_cal1_u143_mac ), .F1(\a_mac_out[6]_cal1_u144_mac ), .F2(\a_mac_out[6]_cal1_u145_mac ), .F3(dummy_abc_369_) );
      defparam ii1190.CONFIG_DATA = 16'h6060;
      defparam ii1190.PLACE_LOCATION = "NONE";
      defparam ii1190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1191 ( .DX(nn1191), .F0(\a_mac_out[6]_cal1_u143_mac ), .F1(\a_mac_out[6]_cal1_u144_mac ), .F2(\a_mac_out[6]_cal1_u145_mac ), .F3(\a_mac_out[6]_cal1_u146_mac ) );
      defparam ii1191.CONFIG_DATA = 16'h9600;
      defparam ii1191.PLACE_LOCATION = "NONE";
      defparam ii1191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1192 ( .DX(nn1192), .F0(\a_mac_out[6]_cal1_u143_mac ), .F1(\a_mac_out[6]_cal1_u144_mac ), .F2(\a_mac_out[7]_cal1_u143_mac ), .F3(\a_mac_out[7]_cal1_u144_mac ) );
      defparam ii1192.CONFIG_DATA = 16'h8778;
      defparam ii1192.PLACE_LOCATION = "NONE";
      defparam ii1192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1193 ( .DX(nn1193), .F0(\a_mac_out[7]_cal1_u145_mac ), .F1(nn1192), .F2(dummy_abc_370_), .F3(dummy_abc_371_) );
      defparam ii1193.CONFIG_DATA = 16'h6666;
      defparam ii1193.PLACE_LOCATION = "NONE";
      defparam ii1193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1194 ( .DX(dOut[1]), .F0(\a_mac_out[7]_cal1_u146_mac ), .F1(nn1190), .F2(nn1191), .F3(nn1193) );
      defparam ii1194.CONFIG_DATA = 16'hA956;
      defparam ii1194.PLACE_LOCATION = "NONE";
      defparam ii1194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1195 ( .DX(nn1195), .F0(\a_mac_out[7]_cal1_u145_mac ), .F1(nn1190), .F2(nn1192), .F3(dummy_abc_372_) );
      defparam ii1195.CONFIG_DATA = 16'hE8E8;
      defparam ii1195.PLACE_LOCATION = "NONE";
      defparam ii1195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1196 ( .DX(nn1196), .F0(\a_mac_out[6]_cal1_u143_mac ), .F1(\a_mac_out[6]_cal1_u144_mac ), .F2(\a_mac_out[7]_cal1_u143_mac ), .F3(\a_mac_out[7]_cal1_u144_mac ) );
      defparam ii1196.CONFIG_DATA = 16'hF880;
      defparam ii1196.PLACE_LOCATION = "NONE";
      defparam ii1196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1197 ( .DX(nn1197), .F0(\a_mac_out[8]_cal1_u143_mac ), .F1(\a_mac_out[8]_cal1_u144_mac ), .F2(\a_mac_out[8]_cal1_u145_mac ), .F3(nn1196) );
      defparam ii1197.CONFIG_DATA = 16'h6996;
      defparam ii1197.PLACE_LOCATION = "NONE";
      defparam ii1197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1198 ( .DX(nn1198), .F0(\a_mac_out[7]_cal1_u146_mac ), .F1(nn1190), .F2(nn1191), .F3(nn1193) );
      defparam ii1198.CONFIG_DATA = 16'hF2A8;
      defparam ii1198.PLACE_LOCATION = "NONE";
      defparam ii1198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1199 ( .DX(dOut[2]), .F0(\a_mac_out[8]_cal1_u146_mac ), .F1(nn1195), .F2(nn1197), .F3(nn1198) );
      defparam ii1199.CONFIG_DATA = 16'h6996;
      defparam ii1199.PLACE_LOCATION = "NONE";
      defparam ii1199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1200 ( .DX(nn1200), .F0(\a_mac_out[8]_cal1_u146_mac ), .F1(nn1195), .F2(nn1197), .F3(nn1198) );
      defparam ii1200.CONFIG_DATA = 16'hBE28;
      defparam ii1200.PLACE_LOCATION = "NONE";
      defparam ii1200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1201 ( .DX(nn1201), .F0(\a_mac_out[8]_cal1_u143_mac ), .F1(\a_mac_out[8]_cal1_u144_mac ), .F2(nn1196), .F3(dummy_abc_373_) );
      defparam ii1201.CONFIG_DATA = 16'hE8E8;
      defparam ii1201.PLACE_LOCATION = "NONE";
      defparam ii1201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1202 ( .DX(nn1202), .F0(\a_mac_out[9]_cal1_u143_mac ), .F1(\a_mac_out[9]_cal1_u144_mac ), .F2(nn1201), .F3(dummy_abc_374_) );
      defparam ii1202.CONFIG_DATA = 16'h6969;
      defparam ii1202.PLACE_LOCATION = "NONE";
      defparam ii1202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1203 ( .DX(nn1203), .F0(\a_mac_out[8]_cal1_u145_mac ), .F1(nn1195), .F2(nn1197), .F3(dummy_abc_375_) );
      defparam ii1203.CONFIG_DATA = 16'h3535;
      defparam ii1203.PLACE_LOCATION = "NONE";
      defparam ii1203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1204 ( .DX(nn1204), .F0(\a_mac_out[9]_cal1_u145_mac ), .F1(nn1202), .F2(nn1203), .F3(dummy_abc_376_) );
      defparam ii1204.CONFIG_DATA = 16'h6969;
      defparam ii1204.PLACE_LOCATION = "NONE";
      defparam ii1204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1205 ( .DX(dOut[3]), .F0(\a_mac_out[9]_cal1_u146_mac ), .F1(nn1200), .F2(nn1204), .F3(dummy_abc_377_) );
      defparam ii1205.CONFIG_DATA = 16'h6969;
      defparam ii1205.PLACE_LOCATION = "NONE";
      defparam ii1205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1206 ( .DX(nn1206), .F0(\a_mac_out[10]_cal1_u143_mac ), .F1(\a_mac_out[10]_cal1_u144_mac ), .F2(\a_mac_out[10]_cal1_u145_mac ), .F3(\a_mac_out[10]_cal1_u146_mac ) );
      defparam ii1206.CONFIG_DATA = 16'h9669;
      defparam ii1206.PLACE_LOCATION = "NONE";
      defparam ii1206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1207 ( .DX(nn1207), .F0(\a_mac_out[9]_cal1_u143_mac ), .F1(\a_mac_out[9]_cal1_u144_mac ), .F2(nn1201), .F3(nn1206) );
      defparam ii1207.CONFIG_DATA = 16'h17E8;
      defparam ii1207.PLACE_LOCATION = "NONE";
      defparam ii1207.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1208 ( .DX(nn1208), .F0(\a_mac_out[9]_cal1_u145_mac ), .F1(nn1202), .F2(nn1203), .F3(nn1207) );
      defparam ii1208.CONFIG_DATA = 16'h2BD4;
      defparam ii1208.PLACE_LOCATION = "NONE";
      defparam ii1208.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1209 ( .DX(dOut[4]), .F0(\a_mac_out[9]_cal1_u146_mac ), .F1(nn1200), .F2(nn1204), .F3(nn1208) );
      defparam ii1209.CONFIG_DATA = 16'h718E;
      defparam ii1209.PLACE_LOCATION = "NONE";
      defparam ii1209.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1210 ( .DX(dOut[5]), .F0(\a_mac_out[6]_cal1_u139_mac ), .F1(\a_mac_out[6]_cal1_u140_mac ), .F2(\a_mac_out[6]_cal1_u141_mac ), .F3(\a_mac_out[6]_cal1_u142_mac ) );
      defparam ii1210.CONFIG_DATA = 16'h6996;
      defparam ii1210.PLACE_LOCATION = "NONE";
      defparam ii1210.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1211 ( .DX(nn1211), .F0(\a_mac_out[6]_cal1_u139_mac ), .F1(\a_mac_out[6]_cal1_u140_mac ), .F2(\a_mac_out[6]_cal1_u141_mac ), .F3(\a_mac_out[6]_cal1_u142_mac ) );
      defparam ii1211.CONFIG_DATA = 16'h9600;
      defparam ii1211.PLACE_LOCATION = "NONE";
      defparam ii1211.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1212 ( .DX(nn1212), .F0(\a_mac_out[6]_cal1_u139_mac ), .F1(\a_mac_out[6]_cal1_u140_mac ), .F2(dummy_abc_378_), .F3(dummy_abc_379_) );
      defparam ii1212.CONFIG_DATA = 16'h8888;
      defparam ii1212.PLACE_LOCATION = "NONE";
      defparam ii1212.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1213 ( .DX(nn1213), .F0(\a_mac_out[6]_cal1_u139_mac ), .F1(\a_mac_out[6]_cal1_u140_mac ), .F2(\a_mac_out[6]_cal1_u141_mac ), .F3(dummy_abc_380_) );
      defparam ii1213.CONFIG_DATA = 16'hE0E0;
      defparam ii1213.PLACE_LOCATION = "NONE";
      defparam ii1213.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1214 ( .DX(nn1214), .F0(\a_mac_out[7]_cal1_u139_mac ), .F1(\a_mac_out[7]_cal1_u140_mac ), .F2(dummy_abc_381_), .F3(dummy_abc_382_) );
      defparam ii1214.CONFIG_DATA = 16'h6666;
      defparam ii1214.PLACE_LOCATION = "NONE";
      defparam ii1214.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1215 ( .DX(nn1215), .F0(\a_mac_out[7]_cal1_u141_mac ), .F1(nn1212), .F2(nn1213), .F3(nn1214) );
      defparam ii1215.CONFIG_DATA = 16'h56A9;
      defparam ii1215.PLACE_LOCATION = "NONE";
      defparam ii1215.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1216 ( .DX(dOut[6]), .F0(\a_mac_out[7]_cal1_u142_mac ), .F1(nn1211), .F2(nn1215), .F3(dummy_abc_383_) );
      defparam ii1216.CONFIG_DATA = 16'h6969;
      defparam ii1216.PLACE_LOCATION = "NONE";
      defparam ii1216.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1217 ( .DX(nn1217), .F0(\a_mac_out[7]_cal1_u142_mac ), .F1(nn1211), .F2(nn1215), .F3(dummy_abc_384_) );
      defparam ii1217.CONFIG_DATA = 16'h7171;
      defparam ii1217.PLACE_LOCATION = "NONE";
      defparam ii1217.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1218 ( .DX(nn1218), .F0(\a_mac_out[7]_cal1_u141_mac ), .F1(nn1212), .F2(nn1213), .F3(nn1214) );
      defparam ii1218.CONFIG_DATA = 16'hCD57;
      defparam ii1218.PLACE_LOCATION = "NONE";
      defparam ii1218.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1219 ( .DX(nn1219), .F0(\a_mac_out[6]_cal1_u139_mac ), .F1(\a_mac_out[6]_cal1_u140_mac ), .F2(\a_mac_out[7]_cal1_u139_mac ), .F3(\a_mac_out[7]_cal1_u140_mac ) );
      defparam ii1219.CONFIG_DATA = 16'hF880;
      defparam ii1219.PLACE_LOCATION = "NONE";
      defparam ii1219.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1220 ( .DX(nn1220), .F0(\a_mac_out[8]_cal1_u139_mac ), .F1(\a_mac_out[8]_cal1_u140_mac ), .F2(nn1218), .F3(nn1219) );
      defparam ii1220.CONFIG_DATA = 16'h9669;
      defparam ii1220.PLACE_LOCATION = "NONE";
      defparam ii1220.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1221 ( .DX(dOut[7]), .F0(\a_mac_out[8]_cal1_u141_mac ), .F1(\a_mac_out[8]_cal1_u142_mac ), .F2(nn1217), .F3(nn1220) );
      defparam ii1221.CONFIG_DATA = 16'h9669;
      defparam ii1221.PLACE_LOCATION = "NONE";
      defparam ii1221.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1222 ( .DX(nn1222), .F0(\a_mac_out[8]_cal1_u139_mac ), .F1(\a_mac_out[8]_cal1_u140_mac ), .F2(dummy_abc_385_), .F3(dummy_abc_386_) );
      defparam ii1222.CONFIG_DATA = 16'h6666;
      defparam ii1222.PLACE_LOCATION = "NONE";
      defparam ii1222.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1223 ( .DX(nn1223), .F0(\a_mac_out[8]_cal1_u141_mac ), .F1(nn1218), .F2(nn1219), .F3(nn1222) );
      defparam ii1223.CONFIG_DATA = 16'hD44D;
      defparam ii1223.PLACE_LOCATION = "NONE";
      defparam ii1223.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1224 ( .DX(nn1224), .F0(\a_mac_out[8]_cal1_u141_mac ), .F1(\a_mac_out[8]_cal1_u142_mac ), .F2(nn1217), .F3(nn1220) );
      defparam ii1224.CONFIG_DATA = 16'hB271;
      defparam ii1224.PLACE_LOCATION = "NONE";
      defparam ii1224.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1225 ( .DX(nn1225), .F0(\a_mac_out[8]_cal1_u139_mac ), .F1(\a_mac_out[8]_cal1_u140_mac ), .F2(nn1219), .F3(dummy_abc_387_) );
      defparam ii1225.CONFIG_DATA = 16'h1717;
      defparam ii1225.PLACE_LOCATION = "NONE";
      defparam ii1225.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1226 ( .DX(nn1226), .F0(\a_mac_out[9]_cal1_u139_mac ), .F1(\a_mac_out[9]_cal1_u140_mac ), .F2(\a_mac_out[9]_cal1_u141_mac ), .F3(nn1225) );
      defparam ii1226.CONFIG_DATA = 16'h9669;
      defparam ii1226.PLACE_LOCATION = "NONE";
      defparam ii1226.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1227 ( .DX(dOut[8]), .F0(\a_mac_out[9]_cal1_u142_mac ), .F1(nn1223), .F2(nn1224), .F3(nn1226) );
      defparam ii1227.CONFIG_DATA = 16'h6996;
      defparam ii1227.PLACE_LOCATION = "NONE";
      defparam ii1227.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1228 ( .DX(nn1228), .F0(\a_mac_out[9]_cal1_u141_mac ), .F1(nn1223), .F2(nn1226), .F3(dummy_abc_388_) );
      defparam ii1228.CONFIG_DATA = 16'hC5C5;
      defparam ii1228.PLACE_LOCATION = "NONE";
      defparam ii1228.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1229 ( .DX(nn1229), .F0(\a_mac_out[9]_cal1_u139_mac ), .F1(\a_mac_out[9]_cal1_u140_mac ), .F2(nn1225), .F3(dummy_abc_389_) );
      defparam ii1229.CONFIG_DATA = 16'h8E8E;
      defparam ii1229.PLACE_LOCATION = "NONE";
      defparam ii1229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1230 ( .DX(nn1230), .F0(\a_mac_out[10]_cal1_u139_mac ), .F1(\a_mac_out[10]_cal1_u140_mac ), .F2(nn1229), .F3(dummy_abc_390_) );
      defparam ii1230.CONFIG_DATA = 16'h9696;
      defparam ii1230.PLACE_LOCATION = "NONE";
      defparam ii1230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1231 ( .DX(nn1231), .F0(\a_mac_out[10]_cal1_u141_mac ), .F1(nn1228), .F2(nn1230), .F3(dummy_abc_391_) );
      defparam ii1231.CONFIG_DATA = 16'h6969;
      defparam ii1231.PLACE_LOCATION = "NONE";
      defparam ii1231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1232 ( .DX(nn1232), .F0(\a_mac_out[9]_cal1_u142_mac ), .F1(nn1223), .F2(nn1224), .F3(nn1226) );
      defparam ii1232.CONFIG_DATA = 16'h8E2B;
      defparam ii1232.PLACE_LOCATION = "NONE";
      defparam ii1232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1233 ( .DX(dOut[9]), .F0(\a_mac_out[10]_cal1_u142_mac ), .F1(nn1231), .F2(nn1232), .F3(dummy_abc_392_) );
      defparam ii1233.CONFIG_DATA = 16'h9696;
      defparam ii1233.PLACE_LOCATION = "NONE";
      defparam ii1233.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1234 ( .DX(nn1234), .F0(\a_mac_out[11]_cal1_u139_mac ), .F1(\a_mac_out[11]_cal1_u140_mac ), .F2(\a_mac_out[11]_cal1_u141_mac ), .F3(\a_mac_out[11]_cal1_u142_mac ) );
      defparam ii1234.CONFIG_DATA = 16'h9669;
      defparam ii1234.PLACE_LOCATION = "NONE";
      defparam ii1234.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1235 ( .DX(nn1235), .F0(\a_mac_out[10]_cal1_u139_mac ), .F1(\a_mac_out[10]_cal1_u140_mac ), .F2(nn1229), .F3(nn1234) );
      defparam ii1235.CONFIG_DATA = 16'hE817;
      defparam ii1235.PLACE_LOCATION = "NONE";
      defparam ii1235.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1236 ( .DX(nn1236), .F0(\a_mac_out[10]_cal1_u141_mac ), .F1(nn1228), .F2(nn1230), .F3(nn1235) );
      defparam ii1236.CONFIG_DATA = 16'h4DB2;
      defparam ii1236.PLACE_LOCATION = "NONE";
      defparam ii1236.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1237 ( .DX(dOut[10]), .F0(\a_mac_out[10]_cal1_u142_mac ), .F1(nn1231), .F2(nn1232), .F3(nn1236) );
      defparam ii1237.CONFIG_DATA = 16'h17E8;
      defparam ii1237.PLACE_LOCATION = "NONE";
      defparam ii1237.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1238 ( .DX(dOut[11]), .F0(\a_mac_out[6]_cal1_u135_mac ), .F1(\a_mac_out[6]_cal1_u136_mac ), .F2(\a_mac_out[6]_cal1_u137_mac ), .F3(\a_mac_out[6]_cal1_u138_mac ) );
      defparam ii1238.CONFIG_DATA = 16'h6996;
      defparam ii1238.PLACE_LOCATION = "NONE";
      defparam ii1238.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1239 ( .DX(nn1239), .F0(\a_mac_out[6]_cal1_u135_mac ), .F1(\a_mac_out[6]_cal1_u136_mac ), .F2(\a_mac_out[6]_cal1_u137_mac ), .F3(\a_mac_out[6]_cal1_u138_mac ) );
      defparam ii1239.CONFIG_DATA = 16'h9600;
      defparam ii1239.PLACE_LOCATION = "NONE";
      defparam ii1239.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1240 ( .DX(nn1240), .F0(\a_mac_out[6]_cal1_u135_mac ), .F1(\a_mac_out[6]_cal1_u136_mac ), .F2(\a_mac_out[6]_cal1_u137_mac ), .F3(dummy_abc_393_) );
      defparam ii1240.CONFIG_DATA = 16'hE8E8;
      defparam ii1240.PLACE_LOCATION = "NONE";
      defparam ii1240.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1241 ( .DX(nn1241), .F0(\a_mac_out[7]_cal1_u135_mac ), .F1(\a_mac_out[7]_cal1_u136_mac ), .F2(\a_mac_out[7]_cal1_u137_mac ), .F3(nn1240) );
      defparam ii1241.CONFIG_DATA = 16'h6996;
      defparam ii1241.PLACE_LOCATION = "NONE";
      defparam ii1241.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1242 ( .DX(dOut[12]), .F0(\a_mac_out[7]_cal1_u138_mac ), .F1(nn1239), .F2(nn1241), .F3(dummy_abc_394_) );
      defparam ii1242.CONFIG_DATA = 16'h9696;
      defparam ii1242.PLACE_LOCATION = "NONE";
      defparam ii1242.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1243 ( .DX(nn1243), .F0(\a_mac_out[7]_cal1_u138_mac ), .F1(nn1239), .F2(nn1241), .F3(dummy_abc_395_) );
      defparam ii1243.CONFIG_DATA = 16'hE8E8;
      defparam ii1243.PLACE_LOCATION = "NONE";
      defparam ii1243.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1244 ( .DX(nn1244), .F0(\a_mac_out[7]_cal1_u135_mac ), .F1(\a_mac_out[7]_cal1_u136_mac ), .F2(dummy_abc_396_), .F3(dummy_abc_397_) );
      defparam ii1244.CONFIG_DATA = 16'h8888;
      defparam ii1244.PLACE_LOCATION = "NONE";
      defparam ii1244.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1245 ( .DX(nn1245), .F0(\a_mac_out[7]_cal1_u135_mac ), .F1(\a_mac_out[7]_cal1_u136_mac ), .F2(\a_mac_out[7]_cal1_u137_mac ), .F3(nn1240) );
      defparam ii1245.CONFIG_DATA = 16'hF660;
      defparam ii1245.PLACE_LOCATION = "NONE";
      defparam ii1245.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1246 ( .DX(nn1246), .F0(\a_mac_out[8]_cal1_u135_mac ), .F1(\a_mac_out[8]_cal1_u136_mac ), .F2(nn1244), .F3(nn1245) );
      defparam ii1246.CONFIG_DATA = 16'h6996;
      defparam ii1246.PLACE_LOCATION = "NONE";
      defparam ii1246.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1247 ( .DX(dOut[13]), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\a_mac_out[8]_cal1_u138_mac ), .F2(nn1243), .F3(nn1246) );
      defparam ii1247.CONFIG_DATA = 16'h6996;
      defparam ii1247.PLACE_LOCATION = "NONE";
      defparam ii1247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1248 ( .DX(nn1248), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\a_mac_out[8]_cal1_u138_mac ), .F2(nn1243), .F3(nn1246) );
      defparam ii1248.CONFIG_DATA = 16'h2B17;
      defparam ii1248.PLACE_LOCATION = "NONE";
      defparam ii1248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1249 ( .DX(nn1249), .F0(\a_mac_out[8]_cal1_u135_mac ), .F1(\a_mac_out[8]_cal1_u136_mac ), .F2(nn1244), .F3(dummy_abc_398_) );
      defparam ii1249.CONFIG_DATA = 16'h9696;
      defparam ii1249.PLACE_LOCATION = "NONE";
      defparam ii1249.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1250 ( .DX(nn1250), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(nn1249), .F2(nn1245), .F3(dummy_abc_399_) );
      defparam ii1250.CONFIG_DATA = 16'hE8E8;
      defparam ii1250.PLACE_LOCATION = "NONE";
      defparam ii1250.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1251 ( .DX(nn1251), .F0(\a_mac_out[7]_cal1_u135_mac ), .F1(\a_mac_out[7]_cal1_u136_mac ), .F2(\a_mac_out[8]_cal1_u135_mac ), .F3(\a_mac_out[8]_cal1_u136_mac ) );
      defparam ii1251.CONFIG_DATA = 16'hF880;
      defparam ii1251.PLACE_LOCATION = "NONE";
      defparam ii1251.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1252 ( .DX(nn1252), .F0(\a_mac_out[9]_cal1_u135_mac ), .F1(\a_mac_out[9]_cal1_u136_mac ), .F2(nn1251), .F3(dummy_abc_400_) );
      defparam ii1252.CONFIG_DATA = 16'h9696;
      defparam ii1252.PLACE_LOCATION = "NONE";
      defparam ii1252.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1253 ( .DX(nn1253), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(nn1250), .F2(nn1252), .F3(dummy_abc_401_) );
      defparam ii1253.CONFIG_DATA = 16'h9696;
      defparam ii1253.PLACE_LOCATION = "NONE";
      defparam ii1253.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1254 ( .DX(dOut[14]), .F0(\a_mac_out[9]_cal1_u138_mac ), .F1(nn1248), .F2(nn1253), .F3(dummy_abc_402_) );
      defparam ii1254.CONFIG_DATA = 16'h6969;
      defparam ii1254.PLACE_LOCATION = "NONE";
      defparam ii1254.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1255 ( .DX(nn1255), .F0(\a_mac_out[10]_cal1_u135_mac ), .F1(\a_mac_out[10]_cal1_u136_mac ), .F2(\a_mac_out[10]_cal1_u137_mac ), .F3(\a_mac_out[10]_cal1_u138_mac ) );
      defparam ii1255.CONFIG_DATA = 16'h9669;
      defparam ii1255.PLACE_LOCATION = "NONE";
      defparam ii1255.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1256 ( .DX(nn1256), .F0(\a_mac_out[9]_cal1_u135_mac ), .F1(\a_mac_out[9]_cal1_u136_mac ), .F2(nn1251), .F3(nn1255) );
      defparam ii1256.CONFIG_DATA = 16'h17E8;
      defparam ii1256.PLACE_LOCATION = "NONE";
      defparam ii1256.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1257 ( .DX(nn1257), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(nn1250), .F2(nn1252), .F3(nn1256) );
      defparam ii1257.CONFIG_DATA = 16'hE817;
      defparam ii1257.PLACE_LOCATION = "NONE";
      defparam ii1257.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1258 ( .DX(dOut[15]), .F0(\a_mac_out[9]_cal1_u138_mac ), .F1(nn1248), .F2(nn1253), .F3(nn1257) );
      defparam ii1258.CONFIG_DATA = 16'h4DB2;
      defparam ii1258.PLACE_LOCATION = "NONE";
      defparam ii1258.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1259 ( .DX(nn1259), .F0(outYRes[0]), .F1(\cal1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_403_), .F3(dummy_abc_404_) );
      defparam ii1259.CONFIG_DATA = 16'h9999;
      defparam ii1259.PLACE_LOCATION = "NONE";
      defparam ii1259.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1260 ( .DX(nn1260), .F0(outYRes[1]), .F1(\cal1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_405_), .F3(dummy_abc_406_) );
      defparam ii1260.CONFIG_DATA = 16'h9999;
      defparam ii1260.PLACE_LOCATION = "NONE";
      defparam ii1260.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1261 ( .DX(nn1261), .F0(outYRes[2]), .F1(\cal1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_407_), .F3(dummy_abc_408_) );
      defparam ii1261.CONFIG_DATA = 16'h9999;
      defparam ii1261.PLACE_LOCATION = "NONE";
      defparam ii1261.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1262 ( .DX(nn1262), .F0(outYRes[3]), .F1(\cal1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_409_), .F3(dummy_abc_410_) );
      defparam ii1262.CONFIG_DATA = 16'h9999;
      defparam ii1262.PLACE_LOCATION = "NONE";
      defparam ii1262.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1263 ( .DX(nn1263), .F0(outYRes[4]), .F1(\cal1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_411_), .F3(dummy_abc_412_) );
      defparam ii1263.CONFIG_DATA = 16'h9999;
      defparam ii1263.PLACE_LOCATION = "NONE";
      defparam ii1263.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1264 ( .DX(nn1264), .F0(outYRes[5]), .F1(\cal1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_413_), .F3(dummy_abc_414_) );
      defparam ii1264.CONFIG_DATA = 16'h9999;
      defparam ii1264.PLACE_LOCATION = "NONE";
      defparam ii1264.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1265 ( .DX(nn1265), .F0(outYRes[6]), .F1(\cal1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_415_), .F3(dummy_abc_416_) );
      defparam ii1265.CONFIG_DATA = 16'h9999;
      defparam ii1265.PLACE_LOCATION = "NONE";
      defparam ii1265.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1266 ( .DX(nn1266), .F0(outYRes[7]), .F1(\cal1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_417_), .F3(dummy_abc_418_) );
      defparam ii1266.CONFIG_DATA = 16'h9999;
      defparam ii1266.PLACE_LOCATION = "NONE";
      defparam ii1266.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1267 ( .DX(nn1267), .F0(outYRes[8]), .F1(\cal1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_419_), .F3(dummy_abc_420_) );
      defparam ii1267.CONFIG_DATA = 16'h9999;
      defparam ii1267.PLACE_LOCATION = "NONE";
      defparam ii1267.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1268 ( .DX(nn1268), .F0(outYRes[9]), .F1(\cal1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_421_), .F3(dummy_abc_422_) );
      defparam ii1268.CONFIG_DATA = 16'h9999;
      defparam ii1268.PLACE_LOCATION = "NONE";
      defparam ii1268.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1269 ( .DX(nn1269), .F0(outYRes[10]), .F1(\cal1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_423_), .F3(dummy_abc_424_) );
      defparam ii1269.CONFIG_DATA = 16'h9999;
      defparam ii1269.PLACE_LOCATION = "NONE";
      defparam ii1269.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1270 ( .DX(nn1270), .F0(dummy_abc_425_), .F1(dummy_abc_426_), .F2(dummy_abc_427_), .F3(dummy_abc_428_) );
      defparam ii1270.CONFIG_DATA = 16'hFFFF;
      defparam ii1270.PLACE_LOCATION = "NONE";
      defparam ii1270.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_6_ ( 
        .CA( {a_acc_en_cal1_u134_mac, outYRes[10], outYRes[9], outYRes[8], 
              outYRes[7], outYRes[6], outYRes[5], outYRes[4], outYRes[3], outYRes[2], 
              outYRes[1], outYRes[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_35_ ), 
        .DX( {nn1270, nn1269, nn1268, nn1267, nn1266, nn1265, nn1264, nn1263, 
              nn1262, nn1261, nn1260, nn1259} ), 
        .SUM( {\cal1_u59_XORCI_11|SUM_net , dummy_36_, dummy_37_, dummy_38_, 
              dummy_39_, dummy_40_, dummy_41_, dummy_42_, dummy_43_, dummy_44_, 
              dummy_45_, dummy_46_} )
      );
    CS_LUT4_PRIM ii1285 ( .DX(nn1285), .F0(outXRes[0]), .F1(\cal1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_429_), .F3(dummy_abc_430_) );
      defparam ii1285.CONFIG_DATA = 16'h9999;
      defparam ii1285.PLACE_LOCATION = "NONE";
      defparam ii1285.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1286 ( .DX(nn1286), .F0(outXRes[1]), .F1(\cal1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_431_), .F3(dummy_abc_432_) );
      defparam ii1286.CONFIG_DATA = 16'h9999;
      defparam ii1286.PLACE_LOCATION = "NONE";
      defparam ii1286.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1287 ( .DX(nn1287), .F0(outXRes[2]), .F1(\cal1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_433_), .F3(dummy_abc_434_) );
      defparam ii1287.CONFIG_DATA = 16'h9999;
      defparam ii1287.PLACE_LOCATION = "NONE";
      defparam ii1287.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1288 ( .DX(nn1288), .F0(outXRes[3]), .F1(\cal1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_435_), .F3(dummy_abc_436_) );
      defparam ii1288.CONFIG_DATA = 16'h9999;
      defparam ii1288.PLACE_LOCATION = "NONE";
      defparam ii1288.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1289 ( .DX(nn1289), .F0(outXRes[4]), .F1(\cal1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_437_), .F3(dummy_abc_438_) );
      defparam ii1289.CONFIG_DATA = 16'h9999;
      defparam ii1289.PLACE_LOCATION = "NONE";
      defparam ii1289.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1290 ( .DX(nn1290), .F0(outXRes[5]), .F1(\cal1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_439_), .F3(dummy_abc_440_) );
      defparam ii1290.CONFIG_DATA = 16'h9999;
      defparam ii1290.PLACE_LOCATION = "NONE";
      defparam ii1290.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1291 ( .DX(nn1291), .F0(outXRes[6]), .F1(\cal1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_441_), .F3(dummy_abc_442_) );
      defparam ii1291.CONFIG_DATA = 16'h9999;
      defparam ii1291.PLACE_LOCATION = "NONE";
      defparam ii1291.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1292 ( .DX(nn1292), .F0(outXRes[7]), .F1(\cal1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_443_), .F3(dummy_abc_444_) );
      defparam ii1292.CONFIG_DATA = 16'h9999;
      defparam ii1292.PLACE_LOCATION = "NONE";
      defparam ii1292.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1293 ( .DX(nn1293), .F0(outXRes[8]), .F1(\cal1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_445_), .F3(dummy_abc_446_) );
      defparam ii1293.CONFIG_DATA = 16'h9999;
      defparam ii1293.PLACE_LOCATION = "NONE";
      defparam ii1293.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1294 ( .DX(nn1294), .F0(outXRes[9]), .F1(\cal1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_447_), .F3(dummy_abc_448_) );
      defparam ii1294.CONFIG_DATA = 16'h9999;
      defparam ii1294.PLACE_LOCATION = "NONE";
      defparam ii1294.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1295 ( .DX(nn1295), .F0(outXRes[10]), .F1(\cal1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_449_), .F3(dummy_abc_450_) );
      defparam ii1295.CONFIG_DATA = 16'h9999;
      defparam ii1295.PLACE_LOCATION = "NONE";
      defparam ii1295.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1296 ( .DX(nn1296), .F0(dummy_abc_451_), .F1(dummy_abc_452_), .F2(dummy_abc_453_), .F3(dummy_abc_454_) );
      defparam ii1296.CONFIG_DATA = 16'hFFFF;
      defparam ii1296.PLACE_LOCATION = "NONE";
      defparam ii1296.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12 ( 
        .CA( {a_acc_en_cal1_u134_mac, outXRes[10], outXRes[9], outXRes[8], 
              outXRes[7], outXRes[6], outXRes[5], outXRes[4], outXRes[3], outXRes[2], 
              outXRes[1], outXRes[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_22_ ), 
        .DX( {nn1296, nn1295, nn1294, nn1293, nn1292, nn1291, nn1290, nn1289, 
              nn1288, nn1287, nn1286, nn1285} ), 
        .SUM( {\cal1_u57_XORCI_11|SUM_net , dummy_23_, dummy_24_, dummy_25_, 
              dummy_26_, dummy_27_, dummy_28_, dummy_29_, dummy_30_, dummy_31_, 
              dummy_32_, dummy_33_} )
      );
    CS_LUT4_PRIM ii1311 ( .DX(nn1311), .F0(HS_1863_net), .F1(\cal1_VSNormal__reg|Q_net ), .F2(\cal1_enforceJmp__reg|Q_net ), .F3(dummy_abc_455_) );
      defparam ii1311.CONFIG_DATA = 16'h0101;
      defparam ii1311.PLACE_LOCATION = "NONE";
      defparam ii1311.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1312 ( .DX(nn1312), .F0(u6810_IN), .F1(dummy_123_), .F2(u3634_OUT), .F3(nn1311) );
      defparam ii1312.CONFIG_DATA = 16'h8F00;
      defparam ii1312.PLACE_LOCATION = "NONE";
      defparam ii1312.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1313 ( .DX(nn1313), .F0(\cal1_xAddress__reg[3]|Q_net ), .F1(\cal1_xAddress__reg[4]|Q_net ), .F2(\cal1_xAddress__reg[5]|Q_net ), .F3(\cal1_xAddress__reg[6]|Q_net ) );
      defparam ii1313.CONFIG_DATA = 16'h0001;
      defparam ii1313.PLACE_LOCATION = "NONE";
      defparam ii1313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1314 ( .DX(nn1314), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(\cal1_xAddress__reg[10]|Q_net ), .F2(\cal1_xAddress__reg[1]|Q_net ), .F3(nn1313) );
      defparam ii1314.CONFIG_DATA = 16'h0100;
      defparam ii1314.PLACE_LOCATION = "NONE";
      defparam ii1314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1315 ( .DX(nn1315), .F0(\cal1_xAddress__reg[7]|Q_net ), .F1(\cal1_xAddress__reg[8]|Q_net ), .F2(\cal1_xAddress__reg[9]|Q_net ), .F3(nn1314) );
      defparam ii1315.CONFIG_DATA = 16'h0100;
      defparam ii1315.PLACE_LOCATION = "NONE";
      defparam ii1315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1316 ( .DX(nn1316), .F0(\cal1_yAddress__reg[3]|Q_net ), .F1(\cal1_yAddress__reg[4]|Q_net ), .F2(\cal1_yAddress__reg[5]|Q_net ), .F3(\cal1_yAddress__reg[6]|Q_net ) );
      defparam ii1316.CONFIG_DATA = 16'h0001;
      defparam ii1316.PLACE_LOCATION = "NONE";
      defparam ii1316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1317 ( .DX(nn1317), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(\cal1_yAddress__reg[10]|Q_net ), .F2(\cal1_yAddress__reg[1]|Q_net ), .F3(nn1316) );
      defparam ii1317.CONFIG_DATA = 16'h0100;
      defparam ii1317.PLACE_LOCATION = "NONE";
      defparam ii1317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1318 ( .DX(nn1318), .F0(\cal1_yAddress__reg[7]|Q_net ), .F1(\cal1_yAddress__reg[8]|Q_net ), .F2(\cal1_yAddress__reg[9]|Q_net ), .F3(nn1317) );
      defparam ii1318.CONFIG_DATA = 16'h0100;
      defparam ii1318.PLACE_LOCATION = "NONE";
      defparam ii1318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1319 ( .DX(nn1319), .F0(\cal1_xAddress__reg[2]|Q_net ), .F1(\cal1_yAddress__reg[2]|Q_net ), .F2(nn1315), .F3(nn1318) );
      defparam ii1319.CONFIG_DATA = 16'h8CAF;
      defparam ii1319.PLACE_LOCATION = "NONE";
      defparam ii1319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1320 ( .DX(dOutEn), .F0(dummy_35_), .F1(dummy_22_), .F2(nn1312), .F3(nn1319) );
      defparam ii1320.CONFIG_DATA = 16'h8000;
      defparam ii1320.PLACE_LOCATION = "NONE";
      defparam ii1320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1321 ( .DX(\haa[0]_fifo1_ram_inst_0_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F2(u6796_O), .F3(nn1092) );
      defparam ii1321.CONFIG_DATA = 16'h00CA;
      defparam ii1321.PLACE_LOCATION = "NONE";
      defparam ii1321.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1322 ( .DX(nn1322), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F2(u3634_OUT), .F3(nn1094) );
      defparam ii1322.CONFIG_DATA = 16'h33F5;
      defparam ii1322.PLACE_LOCATION = "NONE";
      defparam ii1322.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1323 ( .DX(\haa[0]_fifo1_ram_inst_1_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(nn1094), .F2(u3662_O), .F3(nn1322) );
      defparam ii1323.CONFIG_DATA = 16'h20FF;
      defparam ii1323.PLACE_LOCATION = "NONE";
      defparam ii1323.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1324 ( .DX(\haa[0]_fifo1_ram_inst_2_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(nn1094), .F2(u3672_O), .F3(nn1322) );
      defparam ii1324.CONFIG_DATA = 16'h20FF;
      defparam ii1324.PLACE_LOCATION = "NONE";
      defparam ii1324.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1325 ( .DX(u6776_O), .F0(u3634_OUT), .F1(dummy_abc_456_), .F2(dummy_abc_457_), .F3(dummy_abc_458_) );
      defparam ii1325.CONFIG_DATA = 16'h5555;
      defparam ii1325.PLACE_LOCATION = "NONE";
      defparam ii1325.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1326 ( .DX(wea_fifo1_ram_inst_0_u_emb18k_0), .F0(rst), .F1(u4510_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(\inputctrl1_ramWrtEn__reg|Q_net ) );
      defparam ii1326.CONFIG_DATA = 16'hEA00;
      defparam ii1326.PLACE_LOCATION = "NONE";
      defparam ii1326.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1327 ( .DX(wea_fifo1_ram_inst_1_u_emb18k_0), .F0(rst), .F1(u4510_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(\inputctrl1_ramWrtEn__reg|Q_net ) );
      defparam ii1327.CONFIG_DATA = 16'h4000;
      defparam ii1327.PLACE_LOCATION = "NONE";
      defparam ii1327.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1328 ( .DX(nn1328), .F0(dummy_35_), .F1(dummy_22_), .F2(dummy_abc_459_), .F3(dummy_abc_460_) );
      defparam ii1328.CONFIG_DATA = 16'h2222;
      defparam ii1328.PLACE_LOCATION = "NONE";
      defparam ii1328.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1329 ( .DX(nn1329), .F0(dummy_35_), .F1(dummy_22_), .F2(dummy_abc_461_), .F3(dummy_abc_462_) );
      defparam ii1329.CONFIG_DATA = 16'h7777;
      defparam ii1329.PLACE_LOCATION = "NONE";
      defparam ii1329.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1330 ( .DX(nn1330), .F0(\cal1_VSNormal__reg|Q_net ), .F1(dummy_35_), .F2(nn1329), .F3(dummy_abc_463_) );
      defparam ii1330.CONFIG_DATA = 16'hB0B0;
      defparam ii1330.PLACE_LOCATION = "NONE";
      defparam ii1330.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1331 ( .DX(nn1331), .F0(\cal1_jmp1Normal__reg|Q_net ), .F1(dummy_123_), .F2(dummy_abc_464_), .F3(dummy_abc_465_) );
      defparam ii1331.CONFIG_DATA = 16'h1111;
      defparam ii1331.PLACE_LOCATION = "NONE";
      defparam ii1331.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1332 ( .DX(nn1332), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_466_), .F3(dummy_abc_467_) );
      defparam ii1332.CONFIG_DATA = 16'h9999;
      defparam ii1332.PLACE_LOCATION = "NONE";
      defparam ii1332.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1333 ( .DX(nn1333), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_468_), .F3(dummy_abc_469_) );
      defparam ii1333.CONFIG_DATA = 16'h9999;
      defparam ii1333.PLACE_LOCATION = "NONE";
      defparam ii1333.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1334 ( .DX(nn1334), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_abc_470_), .F3(dummy_abc_471_) );
      defparam ii1334.CONFIG_DATA = 16'h9999;
      defparam ii1334.PLACE_LOCATION = "NONE";
      defparam ii1334.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1335 ( .DX(nn1335), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[3]|Q_net ), .F2(dummy_abc_472_), .F3(dummy_abc_473_) );
      defparam ii1335.CONFIG_DATA = 16'h9999;
      defparam ii1335.PLACE_LOCATION = "NONE";
      defparam ii1335.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1336 ( .DX(nn1336), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[4]|Q_net ), .F2(dummy_abc_474_), .F3(dummy_abc_475_) );
      defparam ii1336.CONFIG_DATA = 16'h9999;
      defparam ii1336.PLACE_LOCATION = "NONE";
      defparam ii1336.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1337 ( .DX(nn1337), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[5]|Q_net ), .F2(dummy_abc_476_), .F3(dummy_abc_477_) );
      defparam ii1337.CONFIG_DATA = 16'h9999;
      defparam ii1337.PLACE_LOCATION = "NONE";
      defparam ii1337.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1338 ( .DX(nn1338), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[6]|Q_net ), .F2(dummy_abc_478_), .F3(dummy_abc_479_) );
      defparam ii1338.CONFIG_DATA = 16'h9999;
      defparam ii1338.PLACE_LOCATION = "NONE";
      defparam ii1338.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1339 ( .DX(nn1339), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[7]|Q_net ), .F2(dummy_abc_480_), .F3(dummy_abc_481_) );
      defparam ii1339.CONFIG_DATA = 16'h9999;
      defparam ii1339.PLACE_LOCATION = "NONE";
      defparam ii1339.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1340 ( .DX(nn1340), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[8]|Q_net ), .F2(dummy_abc_482_), .F3(dummy_abc_483_) );
      defparam ii1340.CONFIG_DATA = 16'h9999;
      defparam ii1340.PLACE_LOCATION = "NONE";
      defparam ii1340.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1341 ( .DX(nn1341), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[9]|Q_net ), .F2(dummy_abc_484_), .F3(dummy_abc_485_) );
      defparam ii1341.CONFIG_DATA = 16'h9999;
      defparam ii1341.PLACE_LOCATION = "NONE";
      defparam ii1341.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1342 ( .DX(nn1342), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[10]|Q_net ), .F2(dummy_abc_486_), .F3(dummy_abc_487_) );
      defparam ii1342.CONFIG_DATA = 16'h9999;
      defparam ii1342.PLACE_LOCATION = "NONE";
      defparam ii1342.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1343 ( .DX(nn1343), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[11]|Q_net ), .F2(dummy_abc_488_), .F3(dummy_abc_489_) );
      defparam ii1343.CONFIG_DATA = 16'h9999;
      defparam ii1343.PLACE_LOCATION = "NONE";
      defparam ii1343.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1344 ( .DX(nn1344), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[12]|Q_net ), .F2(dummy_abc_490_), .F3(dummy_abc_491_) );
      defparam ii1344.CONFIG_DATA = 16'h9999;
      defparam ii1344.PLACE_LOCATION = "NONE";
      defparam ii1344.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1345 ( .DX(nn1345), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[13]|Q_net ), .F2(dummy_abc_492_), .F3(dummy_abc_493_) );
      defparam ii1345.CONFIG_DATA = 16'h9999;
      defparam ii1345.PLACE_LOCATION = "NONE";
      defparam ii1345.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1346 ( .DX(nn1346), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[14]|Q_net ), .F2(dummy_abc_494_), .F3(dummy_abc_495_) );
      defparam ii1346.CONFIG_DATA = 16'h9999;
      defparam ii1346.PLACE_LOCATION = "NONE";
      defparam ii1346.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1347 ( .DX(nn1347), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[15]|Q_net ), .F2(dummy_abc_496_), .F3(dummy_abc_497_) );
      defparam ii1347.CONFIG_DATA = 16'h9999;
      defparam ii1347.PLACE_LOCATION = "NONE";
      defparam ii1347.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1348 ( .DX(nn1348), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_498_), .F3(dummy_abc_499_) );
      defparam ii1348.CONFIG_DATA = 16'h9999;
      defparam ii1348.PLACE_LOCATION = "NONE";
      defparam ii1348.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1349 ( .DX(nn1349), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_500_), .F3(dummy_abc_501_) );
      defparam ii1349.CONFIG_DATA = 16'h9999;
      defparam ii1349.PLACE_LOCATION = "NONE";
      defparam ii1349.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1350 ( .DX(nn1350), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_abc_502_), .F2(dummy_abc_503_), .F3(dummy_abc_504_) );
      defparam ii1350.CONFIG_DATA = 16'h5555;
      defparam ii1350.PLACE_LOCATION = "NONE";
      defparam ii1350.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1351 ( .DX(nn1351), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_505_), .F2(dummy_abc_506_), .F3(dummy_abc_507_) );
      defparam ii1351.CONFIG_DATA = 16'h5555;
      defparam ii1351.PLACE_LOCATION = "NONE";
      defparam ii1351.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1352 ( .DX(nn1352), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_508_), .F2(dummy_abc_509_), .F3(dummy_abc_510_) );
      defparam ii1352.CONFIG_DATA = 16'h5555;
      defparam ii1352.PLACE_LOCATION = "NONE";
      defparam ii1352.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1353 ( .DX(nn1353), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_511_), .F2(dummy_abc_512_), .F3(dummy_abc_513_) );
      defparam ii1353.CONFIG_DATA = 16'h5555;
      defparam ii1353.PLACE_LOCATION = "NONE";
      defparam ii1353.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1354 ( .DX(nn1354), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_514_), .F2(dummy_abc_515_), .F3(dummy_abc_516_) );
      defparam ii1354.CONFIG_DATA = 16'h5555;
      defparam ii1354.PLACE_LOCATION = "NONE";
      defparam ii1354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1355 ( .DX(nn1355), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_517_), .F2(dummy_abc_518_), .F3(dummy_abc_519_) );
      defparam ii1355.CONFIG_DATA = 16'h5555;
      defparam ii1355.PLACE_LOCATION = "NONE";
      defparam ii1355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1356 ( .DX(nn1356), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_520_), .F2(dummy_abc_521_), .F3(dummy_abc_522_) );
      defparam ii1356.CONFIG_DATA = 16'h5555;
      defparam ii1356.PLACE_LOCATION = "NONE";
      defparam ii1356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1357 ( .DX(nn1357), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_523_), .F2(dummy_abc_524_), .F3(dummy_abc_525_) );
      defparam ii1357.CONFIG_DATA = 16'h5555;
      defparam ii1357.PLACE_LOCATION = "NONE";
      defparam ii1357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1358 ( .DX(nn1358), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_526_), .F2(dummy_abc_527_), .F3(dummy_abc_528_) );
      defparam ii1358.CONFIG_DATA = 16'h5555;
      defparam ii1358.PLACE_LOCATION = "NONE";
      defparam ii1358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1359 ( .DX(nn1359), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_529_), .F2(dummy_abc_530_), .F3(dummy_abc_531_) );
      defparam ii1359.CONFIG_DATA = 16'h5555;
      defparam ii1359.PLACE_LOCATION = "NONE";
      defparam ii1359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1360 ( .DX(nn1360), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_532_), .F2(dummy_abc_533_), .F3(dummy_abc_534_) );
      defparam ii1360.CONFIG_DATA = 16'h5555;
      defparam ii1360.PLACE_LOCATION = "NONE";
      defparam ii1360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1361 ( .DX(nn1361), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_535_), .F2(dummy_abc_536_), .F3(dummy_abc_537_) );
      defparam ii1361.CONFIG_DATA = 16'h5555;
      defparam ii1361.PLACE_LOCATION = "NONE";
      defparam ii1361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1362 ( .DX(nn1362), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_538_), .F2(dummy_abc_539_), .F3(dummy_abc_540_) );
      defparam ii1362.CONFIG_DATA = 16'h5555;
      defparam ii1362.PLACE_LOCATION = "NONE";
      defparam ii1362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1363 ( .DX(nn1363), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_541_), .F2(dummy_abc_542_), .F3(dummy_abc_543_) );
      defparam ii1363.CONFIG_DATA = 16'h5555;
      defparam ii1363.PLACE_LOCATION = "NONE";
      defparam ii1363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1364 ( .DX(nn1364), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_544_), .F2(dummy_abc_545_), .F3(dummy_abc_546_) );
      defparam ii1364.CONFIG_DATA = 16'h5555;
      defparam ii1364.PLACE_LOCATION = "NONE";
      defparam ii1364.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1365 ( .DX(nn1365), .F0(dummy_abc_547_), .F1(dummy_abc_548_), .F2(dummy_abc_549_), .F3(dummy_abc_550_) );
      defparam ii1365.CONFIG_DATA = 16'hFFFF;
      defparam ii1365.PLACE_LOCATION = "NONE";
      defparam ii1365.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_56_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_545_ ), 
        .DX( {nn1365, nn1364, nn1363, nn1362, nn1361, nn1360, nn1359, nn1358, 
              nn1357, nn1356, nn1355, nn1354, nn1353, nn1352, nn1351, nn1350, 
              nn1349, nn1348} ), 
        .SUM( {\coefcal1_divide_inst2_u120_XORCI_17|SUM_net , dummy_546_, 
              dummy_547_, dummy_548_, dummy_549_, dummy_550_, dummy_551_, dummy_552_, 
              dummy_553_, dummy_554_, dummy_555_, dummy_556_, dummy_557_, dummy_558_, 
              dummy_559_, dummy_560_, dummy_561_, dummy_562_} )
      );
    CS_LUT4_PRIM ii1386 ( .DX(nn1386), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_551_), .F3(dummy_abc_552_) );
      defparam ii1386.CONFIG_DATA = 16'h9999;
      defparam ii1386.PLACE_LOCATION = "NONE";
      defparam ii1386.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1387 ( .DX(nn1387), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_553_), .F3(dummy_abc_554_) );
      defparam ii1387.CONFIG_DATA = 16'h9999;
      defparam ii1387.PLACE_LOCATION = "NONE";
      defparam ii1387.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1388 ( .DX(nn1388), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_abc_555_), .F2(dummy_abc_556_), .F3(dummy_abc_557_) );
      defparam ii1388.CONFIG_DATA = 16'h5555;
      defparam ii1388.PLACE_LOCATION = "NONE";
      defparam ii1388.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1389 ( .DX(nn1389), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_558_), .F2(dummy_abc_559_), .F3(dummy_abc_560_) );
      defparam ii1389.CONFIG_DATA = 16'h5555;
      defparam ii1389.PLACE_LOCATION = "NONE";
      defparam ii1389.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1390 ( .DX(nn1390), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_561_), .F2(dummy_abc_562_), .F3(dummy_abc_563_) );
      defparam ii1390.CONFIG_DATA = 16'h5555;
      defparam ii1390.PLACE_LOCATION = "NONE";
      defparam ii1390.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1391 ( .DX(nn1391), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_564_), .F2(dummy_abc_565_), .F3(dummy_abc_566_) );
      defparam ii1391.CONFIG_DATA = 16'h5555;
      defparam ii1391.PLACE_LOCATION = "NONE";
      defparam ii1391.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1392 ( .DX(nn1392), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_567_), .F2(dummy_abc_568_), .F3(dummy_abc_569_) );
      defparam ii1392.CONFIG_DATA = 16'h5555;
      defparam ii1392.PLACE_LOCATION = "NONE";
      defparam ii1392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1393 ( .DX(nn1393), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_570_), .F2(dummy_abc_571_), .F3(dummy_abc_572_) );
      defparam ii1393.CONFIG_DATA = 16'h5555;
      defparam ii1393.PLACE_LOCATION = "NONE";
      defparam ii1393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1394 ( .DX(nn1394), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_573_), .F2(dummy_abc_574_), .F3(dummy_abc_575_) );
      defparam ii1394.CONFIG_DATA = 16'h5555;
      defparam ii1394.PLACE_LOCATION = "NONE";
      defparam ii1394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1395 ( .DX(nn1395), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_576_), .F2(dummy_abc_577_), .F3(dummy_abc_578_) );
      defparam ii1395.CONFIG_DATA = 16'h5555;
      defparam ii1395.PLACE_LOCATION = "NONE";
      defparam ii1395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1396 ( .DX(nn1396), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_579_), .F2(dummy_abc_580_), .F3(dummy_abc_581_) );
      defparam ii1396.CONFIG_DATA = 16'h5555;
      defparam ii1396.PLACE_LOCATION = "NONE";
      defparam ii1396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1397 ( .DX(nn1397), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_582_), .F2(dummy_abc_583_), .F3(dummy_abc_584_) );
      defparam ii1397.CONFIG_DATA = 16'h5555;
      defparam ii1397.PLACE_LOCATION = "NONE";
      defparam ii1397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1398 ( .DX(nn1398), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_585_), .F2(dummy_abc_586_), .F3(dummy_abc_587_) );
      defparam ii1398.CONFIG_DATA = 16'h5555;
      defparam ii1398.PLACE_LOCATION = "NONE";
      defparam ii1398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1399 ( .DX(nn1399), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_588_), .F2(dummy_abc_589_), .F3(dummy_abc_590_) );
      defparam ii1399.CONFIG_DATA = 16'h5555;
      defparam ii1399.PLACE_LOCATION = "NONE";
      defparam ii1399.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1400 ( .DX(nn1400), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_591_), .F2(dummy_abc_592_), .F3(dummy_abc_593_) );
      defparam ii1400.CONFIG_DATA = 16'h5555;
      defparam ii1400.PLACE_LOCATION = "NONE";
      defparam ii1400.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1401 ( .DX(nn1401), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_594_), .F2(dummy_abc_595_), .F3(dummy_abc_596_) );
      defparam ii1401.CONFIG_DATA = 16'h5555;
      defparam ii1401.PLACE_LOCATION = "NONE";
      defparam ii1401.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1402 ( .DX(nn1402), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_597_), .F2(dummy_abc_598_), .F3(dummy_abc_599_) );
      defparam ii1402.CONFIG_DATA = 16'h5555;
      defparam ii1402.PLACE_LOCATION = "NONE";
      defparam ii1402.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_40_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, \coefcal1_yDividend__reg[16]|Q_net , 
              \coefcal1_yDividend__reg[15]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_168_ ), 
        .DX( {nn1402, nn1401, nn1400, nn1399, nn1398, nn1397, nn1396, nn1395, 
              nn1394, nn1393, nn1392, nn1391, nn1390, nn1389, nn1388, nn1387, 
              nn1386} ), 
        .SUM( {dummy_169_, \coefcal1_divide_inst2_u102_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_14|SUM_net , \coefcal1_divide_inst2_u102_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_12|SUM_net , \coefcal1_divide_inst2_u102_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_10|SUM_net , \coefcal1_divide_inst2_u102_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_8|SUM_net , \coefcal1_divide_inst2_u102_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_6|SUM_net , \coefcal1_divide_inst2_u102_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_4|SUM_net , \coefcal1_divide_inst2_u102_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_2|SUM_net , \coefcal1_divide_inst2_u102_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1422 ( .DX(nn1422), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(dummy_545_), .F2(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ), .F3(dummy_abc_600_) );
      defparam ii1422.CONFIG_DATA = 16'hB8B8;
      defparam ii1422.PLACE_LOCATION = "NONE";
      defparam ii1422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1423 ( .DX(nn1423), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_601_), .F3(dummy_abc_602_) );
      defparam ii1423.CONFIG_DATA = 16'h9999;
      defparam ii1423.PLACE_LOCATION = "NONE";
      defparam ii1423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1424 ( .DX(nn1424), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_545_) );
      defparam ii1424.CONFIG_DATA = 16'hA569;
      defparam ii1424.PLACE_LOCATION = "NONE";
      defparam ii1424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1425 ( .DX(nn1425), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_545_), .F3(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ) );
      defparam ii1425.CONFIG_DATA = 16'h9C93;
      defparam ii1425.PLACE_LOCATION = "NONE";
      defparam ii1425.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1426 ( .DX(nn1426), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_603_), .F2(dummy_abc_604_), .F3(dummy_abc_605_) );
      defparam ii1426.CONFIG_DATA = 16'h5555;
      defparam ii1426.PLACE_LOCATION = "NONE";
      defparam ii1426.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1427 ( .DX(nn1427), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_606_), .F2(dummy_abc_607_), .F3(dummy_abc_608_) );
      defparam ii1427.CONFIG_DATA = 16'h5555;
      defparam ii1427.PLACE_LOCATION = "NONE";
      defparam ii1427.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1428 ( .DX(nn1428), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_609_), .F2(dummy_abc_610_), .F3(dummy_abc_611_) );
      defparam ii1428.CONFIG_DATA = 16'h5555;
      defparam ii1428.PLACE_LOCATION = "NONE";
      defparam ii1428.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1429 ( .DX(nn1429), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_612_), .F2(dummy_abc_613_), .F3(dummy_abc_614_) );
      defparam ii1429.CONFIG_DATA = 16'h5555;
      defparam ii1429.PLACE_LOCATION = "NONE";
      defparam ii1429.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1430 ( .DX(nn1430), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_615_), .F2(dummy_abc_616_), .F3(dummy_abc_617_) );
      defparam ii1430.CONFIG_DATA = 16'h5555;
      defparam ii1430.PLACE_LOCATION = "NONE";
      defparam ii1430.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1431 ( .DX(nn1431), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_618_), .F2(dummy_abc_619_), .F3(dummy_abc_620_) );
      defparam ii1431.CONFIG_DATA = 16'h5555;
      defparam ii1431.PLACE_LOCATION = "NONE";
      defparam ii1431.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1432 ( .DX(nn1432), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_621_), .F2(dummy_abc_622_), .F3(dummy_abc_623_) );
      defparam ii1432.CONFIG_DATA = 16'h5555;
      defparam ii1432.PLACE_LOCATION = "NONE";
      defparam ii1432.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1433 ( .DX(nn1433), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_624_), .F2(dummy_abc_625_), .F3(dummy_abc_626_) );
      defparam ii1433.CONFIG_DATA = 16'h5555;
      defparam ii1433.PLACE_LOCATION = "NONE";
      defparam ii1433.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1434 ( .DX(nn1434), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_627_), .F2(dummy_abc_628_), .F3(dummy_abc_629_) );
      defparam ii1434.CONFIG_DATA = 16'h5555;
      defparam ii1434.PLACE_LOCATION = "NONE";
      defparam ii1434.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1435 ( .DX(nn1435), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_630_), .F2(dummy_abc_631_), .F3(dummy_abc_632_) );
      defparam ii1435.CONFIG_DATA = 16'h5555;
      defparam ii1435.PLACE_LOCATION = "NONE";
      defparam ii1435.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1436 ( .DX(nn1436), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_633_), .F2(dummy_abc_634_), .F3(dummy_abc_635_) );
      defparam ii1436.CONFIG_DATA = 16'h5555;
      defparam ii1436.PLACE_LOCATION = "NONE";
      defparam ii1436.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1437 ( .DX(nn1437), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_636_), .F2(dummy_abc_637_), .F3(dummy_abc_638_) );
      defparam ii1437.CONFIG_DATA = 16'h5555;
      defparam ii1437.PLACE_LOCATION = "NONE";
      defparam ii1437.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1438 ( .DX(nn1438), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_639_), .F2(dummy_abc_640_), .F3(dummy_abc_641_) );
      defparam ii1438.CONFIG_DATA = 16'h5555;
      defparam ii1438.PLACE_LOCATION = "NONE";
      defparam ii1438.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1439 ( .DX(nn1439), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_642_), .F2(dummy_abc_643_), .F3(dummy_abc_644_) );
      defparam ii1439.CONFIG_DATA = 16'h5555;
      defparam ii1439.PLACE_LOCATION = "NONE";
      defparam ii1439.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1440 ( .DX(nn1440), .F0(dummy_abc_645_), .F1(dummy_abc_646_), .F2(dummy_abc_647_), .F3(dummy_abc_648_) );
      defparam ii1440.CONFIG_DATA = 16'hFFFF;
      defparam ii1440.PLACE_LOCATION = "NONE";
      defparam ii1440.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_57_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_564_ ), 
        .DX( {nn1440, nn1439, nn1438, nn1437, nn1436, nn1435, nn1434, nn1433, 
              nn1432, nn1431, nn1430, nn1429, nn1428, nn1427, nn1426, nn1425, 
              nn1424, nn1423} ), 
        .SUM( {\coefcal1_divide_inst2_u122_XORCI_17|SUM_net , dummy_565_, 
              dummy_566_, dummy_567_, dummy_568_, dummy_569_, dummy_570_, dummy_571_, 
              dummy_572_, dummy_573_, dummy_574_, dummy_575_, dummy_576_, dummy_577_, 
              dummy_578_, dummy_579_, dummy_580_, dummy_581_} )
      );
    CS_LUT4_PRIM ii1461 ( .DX(nn1461), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_545_), .F3(dummy_abc_649_) );
      defparam ii1461.CONFIG_DATA = 16'hA6A6;
      defparam ii1461.PLACE_LOCATION = "NONE";
      defparam ii1461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1462 ( .DX(nn1462), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_650_), .F3(dummy_abc_651_) );
      defparam ii1462.CONFIG_DATA = 16'h9999;
      defparam ii1462.PLACE_LOCATION = "NONE";
      defparam ii1462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1463 ( .DX(nn1463), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_545_) );
      defparam ii1463.CONFIG_DATA = 16'hA569;
      defparam ii1463.PLACE_LOCATION = "NONE";
      defparam ii1463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1464 ( .DX(nn1464), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_545_), .F3(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ) );
      defparam ii1464.CONFIG_DATA = 16'h9C93;
      defparam ii1464.PLACE_LOCATION = "NONE";
      defparam ii1464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1465 ( .DX(nn1465), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_652_), .F2(dummy_abc_653_), .F3(dummy_abc_654_) );
      defparam ii1465.CONFIG_DATA = 16'h5555;
      defparam ii1465.PLACE_LOCATION = "NONE";
      defparam ii1465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1466 ( .DX(nn1466), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_655_), .F2(dummy_abc_656_), .F3(dummy_abc_657_) );
      defparam ii1466.CONFIG_DATA = 16'h5555;
      defparam ii1466.PLACE_LOCATION = "NONE";
      defparam ii1466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1467 ( .DX(nn1467), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_658_), .F2(dummy_abc_659_), .F3(dummy_abc_660_) );
      defparam ii1467.CONFIG_DATA = 16'h5555;
      defparam ii1467.PLACE_LOCATION = "NONE";
      defparam ii1467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1468 ( .DX(nn1468), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_661_), .F2(dummy_abc_662_), .F3(dummy_abc_663_) );
      defparam ii1468.CONFIG_DATA = 16'h5555;
      defparam ii1468.PLACE_LOCATION = "NONE";
      defparam ii1468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1469 ( .DX(nn1469), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_664_), .F2(dummy_abc_665_), .F3(dummy_abc_666_) );
      defparam ii1469.CONFIG_DATA = 16'h5555;
      defparam ii1469.PLACE_LOCATION = "NONE";
      defparam ii1469.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1470 ( .DX(nn1470), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_667_), .F2(dummy_abc_668_), .F3(dummy_abc_669_) );
      defparam ii1470.CONFIG_DATA = 16'h5555;
      defparam ii1470.PLACE_LOCATION = "NONE";
      defparam ii1470.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1471 ( .DX(nn1471), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_670_), .F2(dummy_abc_671_), .F3(dummy_abc_672_) );
      defparam ii1471.CONFIG_DATA = 16'h5555;
      defparam ii1471.PLACE_LOCATION = "NONE";
      defparam ii1471.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1472 ( .DX(nn1472), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_673_), .F2(dummy_abc_674_), .F3(dummy_abc_675_) );
      defparam ii1472.CONFIG_DATA = 16'h5555;
      defparam ii1472.PLACE_LOCATION = "NONE";
      defparam ii1472.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1473 ( .DX(nn1473), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_676_), .F2(dummy_abc_677_), .F3(dummy_abc_678_) );
      defparam ii1473.CONFIG_DATA = 16'h5555;
      defparam ii1473.PLACE_LOCATION = "NONE";
      defparam ii1473.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1474 ( .DX(nn1474), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_679_), .F2(dummy_abc_680_), .F3(dummy_abc_681_) );
      defparam ii1474.CONFIG_DATA = 16'h5555;
      defparam ii1474.PLACE_LOCATION = "NONE";
      defparam ii1474.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1475 ( .DX(nn1475), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_682_), .F2(dummy_abc_683_), .F3(dummy_abc_684_) );
      defparam ii1475.CONFIG_DATA = 16'h5555;
      defparam ii1475.PLACE_LOCATION = "NONE";
      defparam ii1475.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1476 ( .DX(nn1476), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_685_), .F2(dummy_abc_686_), .F3(dummy_abc_687_) );
      defparam ii1476.CONFIG_DATA = 16'h5555;
      defparam ii1476.PLACE_LOCATION = "NONE";
      defparam ii1476.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1477 ( .DX(nn1477), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_688_), .F2(dummy_abc_689_), .F3(dummy_abc_690_) );
      defparam ii1477.CONFIG_DATA = 16'h5555;
      defparam ii1477.PLACE_LOCATION = "NONE";
      defparam ii1477.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1478 ( .DX(nn1478), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_691_), .F2(dummy_abc_692_), .F3(dummy_abc_693_) );
      defparam ii1478.CONFIG_DATA = 16'h5555;
      defparam ii1478.PLACE_LOCATION = "NONE";
      defparam ii1478.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_41_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1422, 
              nn1461, \coefcal1_yDividend__reg[14]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_170_ ), 
        .DX( {nn1478, nn1477, nn1476, nn1475, nn1474, nn1473, nn1472, nn1471, 
              nn1470, nn1469, nn1468, nn1467, nn1466, nn1465, nn1464, nn1463, 
              nn1462} ), 
        .SUM( {dummy_171_, \coefcal1_divide_inst2_u103_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_14|SUM_net , \coefcal1_divide_inst2_u103_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_12|SUM_net , \coefcal1_divide_inst2_u103_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_10|SUM_net , \coefcal1_divide_inst2_u103_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_8|SUM_net , \coefcal1_divide_inst2_u103_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_6|SUM_net , \coefcal1_divide_inst2_u103_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_4|SUM_net , \coefcal1_divide_inst2_u103_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_2|SUM_net , \coefcal1_divide_inst2_u103_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1498 ( .DX(nn1498), .F0(nn1422), .F1(dummy_564_), .F2(\coefcal1_divide_inst2_u103_XORCI_2|SUM_net ), .F3(dummy_abc_694_) );
      defparam ii1498.CONFIG_DATA = 16'hB8B8;
      defparam ii1498.PLACE_LOCATION = "NONE";
      defparam ii1498.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1499 ( .DX(nn1499), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_695_), .F3(dummy_abc_696_) );
      defparam ii1499.CONFIG_DATA = 16'h9999;
      defparam ii1499.PLACE_LOCATION = "NONE";
      defparam ii1499.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1500 ( .DX(nn1500), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_564_) );
      defparam ii1500.CONFIG_DATA = 16'hA569;
      defparam ii1500.PLACE_LOCATION = "NONE";
      defparam ii1500.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1501 ( .DX(nn1501), .F0(dummy_564_), .F1(nn1461), .F2(\coefcal1_divide_inst2_u103_XORCI_1|SUM_net ), .F3(dummy_abc_697_) );
      defparam ii1501.CONFIG_DATA = 16'hD8D8;
      defparam ii1501.PLACE_LOCATION = "NONE";
      defparam ii1501.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1502 ( .DX(nn1502), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1501), .F2(dummy_abc_698_), .F3(dummy_abc_699_) );
      defparam ii1502.CONFIG_DATA = 16'h9999;
      defparam ii1502.PLACE_LOCATION = "NONE";
      defparam ii1502.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1503 ( .DX(nn1503), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1498), .F2(dummy_abc_700_), .F3(dummy_abc_701_) );
      defparam ii1503.CONFIG_DATA = 16'h9999;
      defparam ii1503.PLACE_LOCATION = "NONE";
      defparam ii1503.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1504 ( .DX(nn1504), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_702_), .F2(dummy_abc_703_), .F3(dummy_abc_704_) );
      defparam ii1504.CONFIG_DATA = 16'h5555;
      defparam ii1504.PLACE_LOCATION = "NONE";
      defparam ii1504.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1505 ( .DX(nn1505), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_705_), .F2(dummy_abc_706_), .F3(dummy_abc_707_) );
      defparam ii1505.CONFIG_DATA = 16'h5555;
      defparam ii1505.PLACE_LOCATION = "NONE";
      defparam ii1505.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1506 ( .DX(nn1506), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_708_), .F2(dummy_abc_709_), .F3(dummy_abc_710_) );
      defparam ii1506.CONFIG_DATA = 16'h5555;
      defparam ii1506.PLACE_LOCATION = "NONE";
      defparam ii1506.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1507 ( .DX(nn1507), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_711_), .F2(dummy_abc_712_), .F3(dummy_abc_713_) );
      defparam ii1507.CONFIG_DATA = 16'h5555;
      defparam ii1507.PLACE_LOCATION = "NONE";
      defparam ii1507.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1508 ( .DX(nn1508), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_714_), .F2(dummy_abc_715_), .F3(dummy_abc_716_) );
      defparam ii1508.CONFIG_DATA = 16'h5555;
      defparam ii1508.PLACE_LOCATION = "NONE";
      defparam ii1508.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1509 ( .DX(nn1509), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_717_), .F2(dummy_abc_718_), .F3(dummy_abc_719_) );
      defparam ii1509.CONFIG_DATA = 16'h5555;
      defparam ii1509.PLACE_LOCATION = "NONE";
      defparam ii1509.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1510 ( .DX(nn1510), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_720_), .F2(dummy_abc_721_), .F3(dummy_abc_722_) );
      defparam ii1510.CONFIG_DATA = 16'h5555;
      defparam ii1510.PLACE_LOCATION = "NONE";
      defparam ii1510.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1511 ( .DX(nn1511), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_723_), .F2(dummy_abc_724_), .F3(dummy_abc_725_) );
      defparam ii1511.CONFIG_DATA = 16'h5555;
      defparam ii1511.PLACE_LOCATION = "NONE";
      defparam ii1511.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1512 ( .DX(nn1512), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_726_), .F2(dummy_abc_727_), .F3(dummy_abc_728_) );
      defparam ii1512.CONFIG_DATA = 16'h5555;
      defparam ii1512.PLACE_LOCATION = "NONE";
      defparam ii1512.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1513 ( .DX(nn1513), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_729_), .F2(dummy_abc_730_), .F3(dummy_abc_731_) );
      defparam ii1513.CONFIG_DATA = 16'h5555;
      defparam ii1513.PLACE_LOCATION = "NONE";
      defparam ii1513.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1514 ( .DX(nn1514), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_732_), .F2(dummy_abc_733_), .F3(dummy_abc_734_) );
      defparam ii1514.CONFIG_DATA = 16'h5555;
      defparam ii1514.PLACE_LOCATION = "NONE";
      defparam ii1514.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1515 ( .DX(nn1515), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_735_), .F2(dummy_abc_736_), .F3(dummy_abc_737_) );
      defparam ii1515.CONFIG_DATA = 16'h5555;
      defparam ii1515.PLACE_LOCATION = "NONE";
      defparam ii1515.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1516 ( .DX(nn1516), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_738_), .F2(dummy_abc_739_), .F3(dummy_abc_740_) );
      defparam ii1516.CONFIG_DATA = 16'h5555;
      defparam ii1516.PLACE_LOCATION = "NONE";
      defparam ii1516.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1517 ( .DX(nn1517), .F0(dummy_abc_741_), .F1(dummy_abc_742_), .F2(dummy_abc_743_), .F3(dummy_abc_744_) );
      defparam ii1517.CONFIG_DATA = 16'hFFFF;
      defparam ii1517.PLACE_LOCATION = "NONE";
      defparam ii1517.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_58_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_583_ ), 
        .DX( {nn1517, nn1516, nn1515, nn1514, nn1513, nn1512, nn1511, nn1510, 
              nn1509, nn1508, nn1507, nn1506, nn1505, nn1504, nn1503, nn1502, 
              nn1500, nn1499} ), 
        .SUM( {\coefcal1_divide_inst2_u124_XORCI_17|SUM_net , dummy_584_, 
              dummy_585_, dummy_586_, dummy_587_, dummy_588_, dummy_589_, dummy_590_, 
              dummy_591_, dummy_592_, dummy_593_, dummy_594_, dummy_595_, dummy_596_, 
              dummy_597_, dummy_598_, dummy_599_, dummy_600_} )
      );
    CS_LUT4_PRIM ii1538 ( .DX(nn1538), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_564_), .F3(dummy_abc_745_) );
      defparam ii1538.CONFIG_DATA = 16'hA6A6;
      defparam ii1538.PLACE_LOCATION = "NONE";
      defparam ii1538.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1539 ( .DX(nn1539), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_746_), .F3(dummy_abc_747_) );
      defparam ii1539.CONFIG_DATA = 16'h9999;
      defparam ii1539.PLACE_LOCATION = "NONE";
      defparam ii1539.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1540 ( .DX(nn1540), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_564_) );
      defparam ii1540.CONFIG_DATA = 16'hA569;
      defparam ii1540.PLACE_LOCATION = "NONE";
      defparam ii1540.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1541 ( .DX(nn1541), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1501), .F2(dummy_abc_748_), .F3(dummy_abc_749_) );
      defparam ii1541.CONFIG_DATA = 16'h9999;
      defparam ii1541.PLACE_LOCATION = "NONE";
      defparam ii1541.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1542 ( .DX(nn1542), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1498), .F2(dummy_abc_750_), .F3(dummy_abc_751_) );
      defparam ii1542.CONFIG_DATA = 16'h9999;
      defparam ii1542.PLACE_LOCATION = "NONE";
      defparam ii1542.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1543 ( .DX(nn1543), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_752_), .F2(dummy_abc_753_), .F3(dummy_abc_754_) );
      defparam ii1543.CONFIG_DATA = 16'h5555;
      defparam ii1543.PLACE_LOCATION = "NONE";
      defparam ii1543.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1544 ( .DX(nn1544), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_755_), .F2(dummy_abc_756_), .F3(dummy_abc_757_) );
      defparam ii1544.CONFIG_DATA = 16'h5555;
      defparam ii1544.PLACE_LOCATION = "NONE";
      defparam ii1544.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1545 ( .DX(nn1545), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_758_), .F2(dummy_abc_759_), .F3(dummy_abc_760_) );
      defparam ii1545.CONFIG_DATA = 16'h5555;
      defparam ii1545.PLACE_LOCATION = "NONE";
      defparam ii1545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1546 ( .DX(nn1546), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_761_), .F2(dummy_abc_762_), .F3(dummy_abc_763_) );
      defparam ii1546.CONFIG_DATA = 16'h5555;
      defparam ii1546.PLACE_LOCATION = "NONE";
      defparam ii1546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1547 ( .DX(nn1547), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_764_), .F2(dummy_abc_765_), .F3(dummy_abc_766_) );
      defparam ii1547.CONFIG_DATA = 16'h5555;
      defparam ii1547.PLACE_LOCATION = "NONE";
      defparam ii1547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1548 ( .DX(nn1548), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_767_), .F2(dummy_abc_768_), .F3(dummy_abc_769_) );
      defparam ii1548.CONFIG_DATA = 16'h5555;
      defparam ii1548.PLACE_LOCATION = "NONE";
      defparam ii1548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1549 ( .DX(nn1549), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_770_), .F2(dummy_abc_771_), .F3(dummy_abc_772_) );
      defparam ii1549.CONFIG_DATA = 16'h5555;
      defparam ii1549.PLACE_LOCATION = "NONE";
      defparam ii1549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1550 ( .DX(nn1550), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_773_), .F2(dummy_abc_774_), .F3(dummy_abc_775_) );
      defparam ii1550.CONFIG_DATA = 16'h5555;
      defparam ii1550.PLACE_LOCATION = "NONE";
      defparam ii1550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1551 ( .DX(nn1551), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_776_), .F2(dummy_abc_777_), .F3(dummy_abc_778_) );
      defparam ii1551.CONFIG_DATA = 16'h5555;
      defparam ii1551.PLACE_LOCATION = "NONE";
      defparam ii1551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1552 ( .DX(nn1552), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_779_), .F2(dummy_abc_780_), .F3(dummy_abc_781_) );
      defparam ii1552.CONFIG_DATA = 16'h5555;
      defparam ii1552.PLACE_LOCATION = "NONE";
      defparam ii1552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1553 ( .DX(nn1553), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_782_), .F2(dummy_abc_783_), .F3(dummy_abc_784_) );
      defparam ii1553.CONFIG_DATA = 16'h5555;
      defparam ii1553.PLACE_LOCATION = "NONE";
      defparam ii1553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1554 ( .DX(nn1554), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_785_), .F2(dummy_abc_786_), .F3(dummy_abc_787_) );
      defparam ii1554.CONFIG_DATA = 16'h5555;
      defparam ii1554.PLACE_LOCATION = "NONE";
      defparam ii1554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1555 ( .DX(nn1555), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_788_), .F2(dummy_abc_789_), .F3(dummy_abc_790_) );
      defparam ii1555.CONFIG_DATA = 16'h5555;
      defparam ii1555.PLACE_LOCATION = "NONE";
      defparam ii1555.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_42_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1498, nn1501, nn1538, 
              \coefcal1_yDividend__reg[13]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_172_ ), 
        .DX( {nn1555, nn1554, nn1553, nn1552, nn1551, nn1550, nn1549, nn1548, 
              nn1547, nn1546, nn1545, nn1544, nn1543, nn1542, nn1541, nn1540, 
              nn1539} ), 
        .SUM( {dummy_173_, \coefcal1_divide_inst2_u104_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_14|SUM_net , \coefcal1_divide_inst2_u104_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_12|SUM_net , \coefcal1_divide_inst2_u104_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_10|SUM_net , \coefcal1_divide_inst2_u104_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_8|SUM_net , \coefcal1_divide_inst2_u104_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_6|SUM_net , \coefcal1_divide_inst2_u104_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_4|SUM_net , \coefcal1_divide_inst2_u104_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_2|SUM_net , \coefcal1_divide_inst2_u104_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1575 ( .DX(nn1575), .F0(nn1498), .F1(dummy_583_), .F2(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ), .F3(dummy_abc_791_) );
      defparam ii1575.CONFIG_DATA = 16'hB8B8;
      defparam ii1575.PLACE_LOCATION = "NONE";
      defparam ii1575.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1576 ( .DX(nn1576), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_792_), .F3(dummy_abc_793_) );
      defparam ii1576.CONFIG_DATA = 16'h9999;
      defparam ii1576.PLACE_LOCATION = "NONE";
      defparam ii1576.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1577 ( .DX(nn1577), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_583_) );
      defparam ii1577.CONFIG_DATA = 16'hA569;
      defparam ii1577.PLACE_LOCATION = "NONE";
      defparam ii1577.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1578 ( .DX(nn1578), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_583_), .F2(nn1538), .F3(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ) );
      defparam ii1578.CONFIG_DATA = 16'hA695;
      defparam ii1578.PLACE_LOCATION = "NONE";
      defparam ii1578.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1579 ( .DX(nn1579), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1501), .F2(dummy_583_), .F3(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ) );
      defparam ii1579.CONFIG_DATA = 16'h9A95;
      defparam ii1579.PLACE_LOCATION = "NONE";
      defparam ii1579.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1580 ( .DX(nn1580), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1498), .F2(dummy_583_), .F3(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ) );
      defparam ii1580.CONFIG_DATA = 16'h9A95;
      defparam ii1580.PLACE_LOCATION = "NONE";
      defparam ii1580.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1581 ( .DX(nn1581), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_794_), .F2(dummy_abc_795_), .F3(dummy_abc_796_) );
      defparam ii1581.CONFIG_DATA = 16'h5555;
      defparam ii1581.PLACE_LOCATION = "NONE";
      defparam ii1581.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1582 ( .DX(nn1582), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_797_), .F2(dummy_abc_798_), .F3(dummy_abc_799_) );
      defparam ii1582.CONFIG_DATA = 16'h5555;
      defparam ii1582.PLACE_LOCATION = "NONE";
      defparam ii1582.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1583 ( .DX(nn1583), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_800_), .F2(dummy_abc_801_), .F3(dummy_abc_802_) );
      defparam ii1583.CONFIG_DATA = 16'h5555;
      defparam ii1583.PLACE_LOCATION = "NONE";
      defparam ii1583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1584 ( .DX(nn1584), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_803_), .F2(dummy_abc_804_), .F3(dummy_abc_805_) );
      defparam ii1584.CONFIG_DATA = 16'h5555;
      defparam ii1584.PLACE_LOCATION = "NONE";
      defparam ii1584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1585 ( .DX(nn1585), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_806_), .F2(dummy_abc_807_), .F3(dummy_abc_808_) );
      defparam ii1585.CONFIG_DATA = 16'h5555;
      defparam ii1585.PLACE_LOCATION = "NONE";
      defparam ii1585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1586 ( .DX(nn1586), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_809_), .F2(dummy_abc_810_), .F3(dummy_abc_811_) );
      defparam ii1586.CONFIG_DATA = 16'h5555;
      defparam ii1586.PLACE_LOCATION = "NONE";
      defparam ii1586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1587 ( .DX(nn1587), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_812_), .F2(dummy_abc_813_), .F3(dummy_abc_814_) );
      defparam ii1587.CONFIG_DATA = 16'h5555;
      defparam ii1587.PLACE_LOCATION = "NONE";
      defparam ii1587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1588 ( .DX(nn1588), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_815_), .F2(dummy_abc_816_), .F3(dummy_abc_817_) );
      defparam ii1588.CONFIG_DATA = 16'h5555;
      defparam ii1588.PLACE_LOCATION = "NONE";
      defparam ii1588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1589 ( .DX(nn1589), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_818_), .F2(dummy_abc_819_), .F3(dummy_abc_820_) );
      defparam ii1589.CONFIG_DATA = 16'h5555;
      defparam ii1589.PLACE_LOCATION = "NONE";
      defparam ii1589.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1590 ( .DX(nn1590), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_821_), .F2(dummy_abc_822_), .F3(dummy_abc_823_) );
      defparam ii1590.CONFIG_DATA = 16'h5555;
      defparam ii1590.PLACE_LOCATION = "NONE";
      defparam ii1590.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1591 ( .DX(nn1591), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_824_), .F2(dummy_abc_825_), .F3(dummy_abc_826_) );
      defparam ii1591.CONFIG_DATA = 16'h5555;
      defparam ii1591.PLACE_LOCATION = "NONE";
      defparam ii1591.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1592 ( .DX(nn1592), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_827_), .F2(dummy_abc_828_), .F3(dummy_abc_829_) );
      defparam ii1592.CONFIG_DATA = 16'h5555;
      defparam ii1592.PLACE_LOCATION = "NONE";
      defparam ii1592.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1593 ( .DX(nn1593), .F0(dummy_abc_830_), .F1(dummy_abc_831_), .F2(dummy_abc_832_), .F3(dummy_abc_833_) );
      defparam ii1593.CONFIG_DATA = 16'hFFFF;
      defparam ii1593.PLACE_LOCATION = "NONE";
      defparam ii1593.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_59_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_602_ ), 
        .DX( {nn1593, nn1592, nn1591, nn1590, nn1589, nn1588, nn1587, nn1586, 
              nn1585, nn1584, nn1583, nn1582, nn1581, nn1580, nn1579, nn1578, 
              nn1577, nn1576} ), 
        .SUM( {\coefcal1_divide_inst2_u126_XORCI_17|SUM_net , dummy_603_, 
              dummy_604_, dummy_605_, dummy_606_, dummy_607_, dummy_608_, dummy_609_, 
              dummy_610_, dummy_611_, dummy_612_, dummy_613_, dummy_614_, dummy_615_, 
              dummy_616_, dummy_617_, dummy_618_, dummy_619_} )
      );
    CS_LUT4_PRIM ii1614 ( .DX(nn1614), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_583_), .F3(dummy_abc_834_) );
      defparam ii1614.CONFIG_DATA = 16'hA6A6;
      defparam ii1614.PLACE_LOCATION = "NONE";
      defparam ii1614.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1615 ( .DX(nn1615), .F0(dummy_583_), .F1(nn1538), .F2(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ), .F3(dummy_abc_835_) );
      defparam ii1615.CONFIG_DATA = 16'hD8D8;
      defparam ii1615.PLACE_LOCATION = "NONE";
      defparam ii1615.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1616 ( .DX(nn1616), .F0(nn1501), .F1(dummy_583_), .F2(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ), .F3(dummy_abc_836_) );
      defparam ii1616.CONFIG_DATA = 16'hB8B8;
      defparam ii1616.PLACE_LOCATION = "NONE";
      defparam ii1616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1617 ( .DX(nn1617), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_837_), .F3(dummy_abc_838_) );
      defparam ii1617.CONFIG_DATA = 16'h9999;
      defparam ii1617.PLACE_LOCATION = "NONE";
      defparam ii1617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1618 ( .DX(nn1618), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_583_) );
      defparam ii1618.CONFIG_DATA = 16'hA569;
      defparam ii1618.PLACE_LOCATION = "NONE";
      defparam ii1618.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1619 ( .DX(nn1619), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_583_), .F2(nn1538), .F3(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ) );
      defparam ii1619.CONFIG_DATA = 16'hA695;
      defparam ii1619.PLACE_LOCATION = "NONE";
      defparam ii1619.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1620 ( .DX(nn1620), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1501), .F2(dummy_583_), .F3(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ) );
      defparam ii1620.CONFIG_DATA = 16'h9A95;
      defparam ii1620.PLACE_LOCATION = "NONE";
      defparam ii1620.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1621 ( .DX(nn1621), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1498), .F2(dummy_583_), .F3(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ) );
      defparam ii1621.CONFIG_DATA = 16'h9A95;
      defparam ii1621.PLACE_LOCATION = "NONE";
      defparam ii1621.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1622 ( .DX(nn1622), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_839_), .F2(dummy_abc_840_), .F3(dummy_abc_841_) );
      defparam ii1622.CONFIG_DATA = 16'h5555;
      defparam ii1622.PLACE_LOCATION = "NONE";
      defparam ii1622.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1623 ( .DX(nn1623), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_842_), .F2(dummy_abc_843_), .F3(dummy_abc_844_) );
      defparam ii1623.CONFIG_DATA = 16'h5555;
      defparam ii1623.PLACE_LOCATION = "NONE";
      defparam ii1623.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1624 ( .DX(nn1624), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_845_), .F2(dummy_abc_846_), .F3(dummy_abc_847_) );
      defparam ii1624.CONFIG_DATA = 16'h5555;
      defparam ii1624.PLACE_LOCATION = "NONE";
      defparam ii1624.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1625 ( .DX(nn1625), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_848_), .F2(dummy_abc_849_), .F3(dummy_abc_850_) );
      defparam ii1625.CONFIG_DATA = 16'h5555;
      defparam ii1625.PLACE_LOCATION = "NONE";
      defparam ii1625.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1626 ( .DX(nn1626), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_851_), .F2(dummy_abc_852_), .F3(dummy_abc_853_) );
      defparam ii1626.CONFIG_DATA = 16'h5555;
      defparam ii1626.PLACE_LOCATION = "NONE";
      defparam ii1626.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1627 ( .DX(nn1627), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_854_), .F2(dummy_abc_855_), .F3(dummy_abc_856_) );
      defparam ii1627.CONFIG_DATA = 16'h5555;
      defparam ii1627.PLACE_LOCATION = "NONE";
      defparam ii1627.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1628 ( .DX(nn1628), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_857_), .F2(dummy_abc_858_), .F3(dummy_abc_859_) );
      defparam ii1628.CONFIG_DATA = 16'h5555;
      defparam ii1628.PLACE_LOCATION = "NONE";
      defparam ii1628.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1629 ( .DX(nn1629), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_860_), .F2(dummy_abc_861_), .F3(dummy_abc_862_) );
      defparam ii1629.CONFIG_DATA = 16'h5555;
      defparam ii1629.PLACE_LOCATION = "NONE";
      defparam ii1629.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1630 ( .DX(nn1630), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_863_), .F2(dummy_abc_864_), .F3(dummy_abc_865_) );
      defparam ii1630.CONFIG_DATA = 16'h5555;
      defparam ii1630.PLACE_LOCATION = "NONE";
      defparam ii1630.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1631 ( .DX(nn1631), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_866_), .F2(dummy_abc_867_), .F3(dummy_abc_868_) );
      defparam ii1631.CONFIG_DATA = 16'h5555;
      defparam ii1631.PLACE_LOCATION = "NONE";
      defparam ii1631.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1632 ( .DX(nn1632), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_869_), .F2(dummy_abc_870_), .F3(dummy_abc_871_) );
      defparam ii1632.CONFIG_DATA = 16'h5555;
      defparam ii1632.PLACE_LOCATION = "NONE";
      defparam ii1632.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1633 ( .DX(nn1633), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_872_), .F2(dummy_abc_873_), .F3(dummy_abc_874_) );
      defparam ii1633.CONFIG_DATA = 16'h5555;
      defparam ii1633.PLACE_LOCATION = "NONE";
      defparam ii1633.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_43_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn1575, nn1616, nn1615, nn1614, 
              \coefcal1_yDividend__reg[12]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_174_ ), 
        .DX( {nn1633, nn1632, nn1631, nn1630, nn1629, nn1628, nn1627, nn1626, 
              nn1625, nn1624, nn1623, nn1622, nn1621, nn1620, nn1619, nn1618, 
              nn1617} ), 
        .SUM( {dummy_175_, \coefcal1_divide_inst2_u105_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_14|SUM_net , \coefcal1_divide_inst2_u105_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_12|SUM_net , \coefcal1_divide_inst2_u105_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_10|SUM_net , \coefcal1_divide_inst2_u105_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_8|SUM_net , \coefcal1_divide_inst2_u105_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_6|SUM_net , \coefcal1_divide_inst2_u105_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_4|SUM_net , \coefcal1_divide_inst2_u105_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_2|SUM_net , \coefcal1_divide_inst2_u105_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1653 ( .DX(nn1653), .F0(dummy_602_), .F1(\coefcal1_divide_inst2_u105_XORCI_4|SUM_net ), .F2(dummy_abc_875_), .F3(dummy_abc_876_) );
      defparam ii1653.CONFIG_DATA = 16'h1111;
      defparam ii1653.PLACE_LOCATION = "NONE";
      defparam ii1653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1654 ( .DX(nn1654), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_877_), .F3(dummy_abc_878_) );
      defparam ii1654.CONFIG_DATA = 16'h9999;
      defparam ii1654.PLACE_LOCATION = "NONE";
      defparam ii1654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1655 ( .DX(nn1655), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_602_) );
      defparam ii1655.CONFIG_DATA = 16'hA569;
      defparam ii1655.PLACE_LOCATION = "NONE";
      defparam ii1655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1656 ( .DX(nn1656), .F0(dummy_602_), .F1(nn1614), .F2(\coefcal1_divide_inst2_u105_XORCI_1|SUM_net ), .F3(dummy_abc_879_) );
      defparam ii1656.CONFIG_DATA = 16'hD8D8;
      defparam ii1656.PLACE_LOCATION = "NONE";
      defparam ii1656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1657 ( .DX(nn1657), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1656), .F2(dummy_abc_880_), .F3(dummy_abc_881_) );
      defparam ii1657.CONFIG_DATA = 16'h9999;
      defparam ii1657.PLACE_LOCATION = "NONE";
      defparam ii1657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1658 ( .DX(nn1658), .F0(nn1615), .F1(dummy_602_), .F2(\coefcal1_divide_inst2_u105_XORCI_2|SUM_net ), .F3(dummy_abc_882_) );
      defparam ii1658.CONFIG_DATA = 16'hB8B8;
      defparam ii1658.PLACE_LOCATION = "NONE";
      defparam ii1658.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1659 ( .DX(nn1659), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1658), .F2(dummy_abc_883_), .F3(dummy_abc_884_) );
      defparam ii1659.CONFIG_DATA = 16'h9999;
      defparam ii1659.PLACE_LOCATION = "NONE";
      defparam ii1659.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1660 ( .DX(nn1660), .F0(nn1616), .F1(dummy_602_), .F2(\coefcal1_divide_inst2_u105_XORCI_3|SUM_net ), .F3(dummy_abc_885_) );
      defparam ii1660.CONFIG_DATA = 16'hB8B8;
      defparam ii1660.PLACE_LOCATION = "NONE";
      defparam ii1660.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1661 ( .DX(nn1661), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1660), .F2(dummy_abc_886_), .F3(dummy_abc_887_) );
      defparam ii1661.CONFIG_DATA = 16'h9999;
      defparam ii1661.PLACE_LOCATION = "NONE";
      defparam ii1661.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1662 ( .DX(nn1662), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1575), .F2(nn1653), .F3(dummy_abc_888_) );
      defparam ii1662.CONFIG_DATA = 16'hD9D9;
      defparam ii1662.PLACE_LOCATION = "NONE";
      defparam ii1662.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1663 ( .DX(nn1663), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_889_), .F2(dummy_abc_890_), .F3(dummy_abc_891_) );
      defparam ii1663.CONFIG_DATA = 16'h5555;
      defparam ii1663.PLACE_LOCATION = "NONE";
      defparam ii1663.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1664 ( .DX(nn1664), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_892_), .F2(dummy_abc_893_), .F3(dummy_abc_894_) );
      defparam ii1664.CONFIG_DATA = 16'h5555;
      defparam ii1664.PLACE_LOCATION = "NONE";
      defparam ii1664.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1665 ( .DX(nn1665), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_895_), .F2(dummy_abc_896_), .F3(dummy_abc_897_) );
      defparam ii1665.CONFIG_DATA = 16'h5555;
      defparam ii1665.PLACE_LOCATION = "NONE";
      defparam ii1665.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1666 ( .DX(nn1666), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_898_), .F2(dummy_abc_899_), .F3(dummy_abc_900_) );
      defparam ii1666.CONFIG_DATA = 16'h5555;
      defparam ii1666.PLACE_LOCATION = "NONE";
      defparam ii1666.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1667 ( .DX(nn1667), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_901_), .F2(dummy_abc_902_), .F3(dummy_abc_903_) );
      defparam ii1667.CONFIG_DATA = 16'h5555;
      defparam ii1667.PLACE_LOCATION = "NONE";
      defparam ii1667.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1668 ( .DX(nn1668), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_904_), .F2(dummy_abc_905_), .F3(dummy_abc_906_) );
      defparam ii1668.CONFIG_DATA = 16'h5555;
      defparam ii1668.PLACE_LOCATION = "NONE";
      defparam ii1668.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1669 ( .DX(nn1669), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_907_), .F2(dummy_abc_908_), .F3(dummy_abc_909_) );
      defparam ii1669.CONFIG_DATA = 16'h5555;
      defparam ii1669.PLACE_LOCATION = "NONE";
      defparam ii1669.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1670 ( .DX(nn1670), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_910_), .F2(dummy_abc_911_), .F3(dummy_abc_912_) );
      defparam ii1670.CONFIG_DATA = 16'h5555;
      defparam ii1670.PLACE_LOCATION = "NONE";
      defparam ii1670.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1671 ( .DX(nn1671), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_913_), .F2(dummy_abc_914_), .F3(dummy_abc_915_) );
      defparam ii1671.CONFIG_DATA = 16'h5555;
      defparam ii1671.PLACE_LOCATION = "NONE";
      defparam ii1671.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1672 ( .DX(nn1672), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_916_), .F2(dummy_abc_917_), .F3(dummy_abc_918_) );
      defparam ii1672.CONFIG_DATA = 16'h5555;
      defparam ii1672.PLACE_LOCATION = "NONE";
      defparam ii1672.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1673 ( .DX(nn1673), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_919_), .F2(dummy_abc_920_), .F3(dummy_abc_921_) );
      defparam ii1673.CONFIG_DATA = 16'h5555;
      defparam ii1673.PLACE_LOCATION = "NONE";
      defparam ii1673.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1674 ( .DX(nn1674), .F0(dummy_abc_922_), .F1(dummy_abc_923_), .F2(dummy_abc_924_), .F3(dummy_abc_925_) );
      defparam ii1674.CONFIG_DATA = 16'hFFFF;
      defparam ii1674.PLACE_LOCATION = "NONE";
      defparam ii1674.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_60_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_621_ ), 
        .DX( {nn1674, nn1673, nn1672, nn1671, nn1670, nn1669, nn1668, nn1667, 
              nn1666, nn1665, nn1664, nn1663, nn1662, nn1661, nn1659, nn1657, 
              nn1655, nn1654} ), 
        .SUM( {\coefcal1_divide_inst2_u128_XORCI_17|SUM_net , dummy_622_, 
              dummy_623_, dummy_624_, dummy_625_, dummy_626_, dummy_627_, dummy_628_, 
              dummy_629_, dummy_630_, dummy_631_, dummy_632_, dummy_633_, dummy_634_, 
              dummy_635_, dummy_636_, dummy_637_, dummy_638_} )
      );
    CS_LUT4_PRIM ii1695 ( .DX(nn1695), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_602_), .F3(dummy_abc_926_) );
      defparam ii1695.CONFIG_DATA = 16'hA6A6;
      defparam ii1695.PLACE_LOCATION = "NONE";
      defparam ii1695.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1696 ( .DX(nn1696), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_927_), .F3(dummy_abc_928_) );
      defparam ii1696.CONFIG_DATA = 16'h9999;
      defparam ii1696.PLACE_LOCATION = "NONE";
      defparam ii1696.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1697 ( .DX(nn1697), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_602_) );
      defparam ii1697.CONFIG_DATA = 16'hA569;
      defparam ii1697.PLACE_LOCATION = "NONE";
      defparam ii1697.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1698 ( .DX(nn1698), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1656), .F2(dummy_abc_929_), .F3(dummy_abc_930_) );
      defparam ii1698.CONFIG_DATA = 16'h9999;
      defparam ii1698.PLACE_LOCATION = "NONE";
      defparam ii1698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1699 ( .DX(nn1699), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1658), .F2(dummy_abc_931_), .F3(dummy_abc_932_) );
      defparam ii1699.CONFIG_DATA = 16'h9999;
      defparam ii1699.PLACE_LOCATION = "NONE";
      defparam ii1699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1700 ( .DX(nn1700), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1660), .F2(dummy_abc_933_), .F3(dummy_abc_934_) );
      defparam ii1700.CONFIG_DATA = 16'h9999;
      defparam ii1700.PLACE_LOCATION = "NONE";
      defparam ii1700.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1701 ( .DX(nn1701), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1575), .F2(nn1653), .F3(dummy_abc_935_) );
      defparam ii1701.CONFIG_DATA = 16'hD9D9;
      defparam ii1701.PLACE_LOCATION = "NONE";
      defparam ii1701.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1702 ( .DX(nn1702), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_936_), .F2(dummy_abc_937_), .F3(dummy_abc_938_) );
      defparam ii1702.CONFIG_DATA = 16'h5555;
      defparam ii1702.PLACE_LOCATION = "NONE";
      defparam ii1702.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1703 ( .DX(nn1703), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_939_), .F2(dummy_abc_940_), .F3(dummy_abc_941_) );
      defparam ii1703.CONFIG_DATA = 16'h5555;
      defparam ii1703.PLACE_LOCATION = "NONE";
      defparam ii1703.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1704 ( .DX(nn1704), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_942_), .F2(dummy_abc_943_), .F3(dummy_abc_944_) );
      defparam ii1704.CONFIG_DATA = 16'h5555;
      defparam ii1704.PLACE_LOCATION = "NONE";
      defparam ii1704.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1705 ( .DX(nn1705), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_945_), .F2(dummy_abc_946_), .F3(dummy_abc_947_) );
      defparam ii1705.CONFIG_DATA = 16'h5555;
      defparam ii1705.PLACE_LOCATION = "NONE";
      defparam ii1705.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1706 ( .DX(nn1706), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_948_), .F2(dummy_abc_949_), .F3(dummy_abc_950_) );
      defparam ii1706.CONFIG_DATA = 16'h5555;
      defparam ii1706.PLACE_LOCATION = "NONE";
      defparam ii1706.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1707 ( .DX(nn1707), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_951_), .F2(dummy_abc_952_), .F3(dummy_abc_953_) );
      defparam ii1707.CONFIG_DATA = 16'h5555;
      defparam ii1707.PLACE_LOCATION = "NONE";
      defparam ii1707.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1708 ( .DX(nn1708), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_954_), .F2(dummy_abc_955_), .F3(dummy_abc_956_) );
      defparam ii1708.CONFIG_DATA = 16'h5555;
      defparam ii1708.PLACE_LOCATION = "NONE";
      defparam ii1708.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1709 ( .DX(nn1709), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_957_), .F2(dummy_abc_958_), .F3(dummy_abc_959_) );
      defparam ii1709.CONFIG_DATA = 16'h5555;
      defparam ii1709.PLACE_LOCATION = "NONE";
      defparam ii1709.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1710 ( .DX(nn1710), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_960_), .F2(dummy_abc_961_), .F3(dummy_abc_962_) );
      defparam ii1710.CONFIG_DATA = 16'h5555;
      defparam ii1710.PLACE_LOCATION = "NONE";
      defparam ii1710.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1711 ( .DX(nn1711), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_963_), .F2(dummy_abc_964_), .F3(dummy_abc_965_) );
      defparam ii1711.CONFIG_DATA = 16'h5555;
      defparam ii1711.PLACE_LOCATION = "NONE";
      defparam ii1711.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1712 ( .DX(nn1712), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_966_), .F2(dummy_abc_967_), .F3(dummy_abc_968_) );
      defparam ii1712.CONFIG_DATA = 16'h5555;
      defparam ii1712.PLACE_LOCATION = "NONE";
      defparam ii1712.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_44_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn1660, nn1658, nn1656, nn1695, 
              \coefcal1_yDividend__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_176_ ), 
        .DX( {nn1712, nn1711, nn1710, nn1709, nn1708, nn1707, nn1706, nn1705, 
              nn1704, nn1703, nn1702, nn1701, nn1700, nn1699, nn1698, nn1697, 
              nn1696} ), 
        .SUM( {dummy_177_, \coefcal1_divide_inst2_u106_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_14|SUM_net , \coefcal1_divide_inst2_u106_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_12|SUM_net , \coefcal1_divide_inst2_u106_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_10|SUM_net , \coefcal1_divide_inst2_u106_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_8|SUM_net , \coefcal1_divide_inst2_u106_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_6|SUM_net , \coefcal1_divide_inst2_u106_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_4|SUM_net , \coefcal1_divide_inst2_u106_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_2|SUM_net , \coefcal1_divide_inst2_u106_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1732 ( .DX(nn1732), .F0(nn1575), .F1(nn1653), .F2(dummy_621_), .F3(\coefcal1_divide_inst2_u106_XORCI_5|SUM_net ) );
      defparam ii1732.CONFIG_DATA = 16'h2A20;
      defparam ii1732.PLACE_LOCATION = "NONE";
      defparam ii1732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1733 ( .DX(nn1733), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_969_), .F3(dummy_abc_970_) );
      defparam ii1733.CONFIG_DATA = 16'h9999;
      defparam ii1733.PLACE_LOCATION = "NONE";
      defparam ii1733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1734 ( .DX(nn1734), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_621_) );
      defparam ii1734.CONFIG_DATA = 16'hA569;
      defparam ii1734.PLACE_LOCATION = "NONE";
      defparam ii1734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1735 ( .DX(nn1735), .F0(dummy_621_), .F1(nn1695), .F2(\coefcal1_divide_inst2_u106_XORCI_1|SUM_net ), .F3(dummy_abc_971_) );
      defparam ii1735.CONFIG_DATA = 16'hD8D8;
      defparam ii1735.PLACE_LOCATION = "NONE";
      defparam ii1735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1736 ( .DX(nn1736), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1735), .F2(dummy_abc_972_), .F3(dummy_abc_973_) );
      defparam ii1736.CONFIG_DATA = 16'h9999;
      defparam ii1736.PLACE_LOCATION = "NONE";
      defparam ii1736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1737 ( .DX(nn1737), .F0(nn1656), .F1(dummy_621_), .F2(\coefcal1_divide_inst2_u106_XORCI_2|SUM_net ), .F3(dummy_abc_974_) );
      defparam ii1737.CONFIG_DATA = 16'hB8B8;
      defparam ii1737.PLACE_LOCATION = "NONE";
      defparam ii1737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1738 ( .DX(nn1738), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1737), .F2(dummy_abc_975_), .F3(dummy_abc_976_) );
      defparam ii1738.CONFIG_DATA = 16'h9999;
      defparam ii1738.PLACE_LOCATION = "NONE";
      defparam ii1738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1739 ( .DX(nn1739), .F0(nn1658), .F1(dummy_621_), .F2(\coefcal1_divide_inst2_u106_XORCI_3|SUM_net ), .F3(dummy_abc_977_) );
      defparam ii1739.CONFIG_DATA = 16'hB8B8;
      defparam ii1739.PLACE_LOCATION = "NONE";
      defparam ii1739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1740 ( .DX(nn1740), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1739), .F2(dummy_abc_978_), .F3(dummy_abc_979_) );
      defparam ii1740.CONFIG_DATA = 16'h9999;
      defparam ii1740.PLACE_LOCATION = "NONE";
      defparam ii1740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1741 ( .DX(nn1741), .F0(nn1660), .F1(dummy_621_), .F2(\coefcal1_divide_inst2_u106_XORCI_4|SUM_net ), .F3(dummy_abc_980_) );
      defparam ii1741.CONFIG_DATA = 16'hB8B8;
      defparam ii1741.PLACE_LOCATION = "NONE";
      defparam ii1741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1742 ( .DX(nn1742), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1741), .F2(dummy_abc_981_), .F3(dummy_abc_982_) );
      defparam ii1742.CONFIG_DATA = 16'h9999;
      defparam ii1742.PLACE_LOCATION = "NONE";
      defparam ii1742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1743 ( .DX(nn1743), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1732), .F2(dummy_abc_983_), .F3(dummy_abc_984_) );
      defparam ii1743.CONFIG_DATA = 16'h9999;
      defparam ii1743.PLACE_LOCATION = "NONE";
      defparam ii1743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1744 ( .DX(nn1744), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_985_), .F2(dummy_abc_986_), .F3(dummy_abc_987_) );
      defparam ii1744.CONFIG_DATA = 16'h5555;
      defparam ii1744.PLACE_LOCATION = "NONE";
      defparam ii1744.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1745 ( .DX(nn1745), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_988_), .F2(dummy_abc_989_), .F3(dummy_abc_990_) );
      defparam ii1745.CONFIG_DATA = 16'h5555;
      defparam ii1745.PLACE_LOCATION = "NONE";
      defparam ii1745.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1746 ( .DX(nn1746), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_991_), .F2(dummy_abc_992_), .F3(dummy_abc_993_) );
      defparam ii1746.CONFIG_DATA = 16'h5555;
      defparam ii1746.PLACE_LOCATION = "NONE";
      defparam ii1746.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1747 ( .DX(nn1747), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_994_), .F2(dummy_abc_995_), .F3(dummy_abc_996_) );
      defparam ii1747.CONFIG_DATA = 16'h5555;
      defparam ii1747.PLACE_LOCATION = "NONE";
      defparam ii1747.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1748 ( .DX(nn1748), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_997_), .F2(dummy_abc_998_), .F3(dummy_abc_999_) );
      defparam ii1748.CONFIG_DATA = 16'h5555;
      defparam ii1748.PLACE_LOCATION = "NONE";
      defparam ii1748.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1749 ( .DX(nn1749), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1000_), .F2(dummy_abc_1001_), .F3(dummy_abc_1002_) );
      defparam ii1749.CONFIG_DATA = 16'h5555;
      defparam ii1749.PLACE_LOCATION = "NONE";
      defparam ii1749.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1750 ( .DX(nn1750), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1003_), .F2(dummy_abc_1004_), .F3(dummy_abc_1005_) );
      defparam ii1750.CONFIG_DATA = 16'h5555;
      defparam ii1750.PLACE_LOCATION = "NONE";
      defparam ii1750.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1751 ( .DX(nn1751), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1006_), .F2(dummy_abc_1007_), .F3(dummy_abc_1008_) );
      defparam ii1751.CONFIG_DATA = 16'h5555;
      defparam ii1751.PLACE_LOCATION = "NONE";
      defparam ii1751.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1752 ( .DX(nn1752), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1009_), .F2(dummy_abc_1010_), .F3(dummy_abc_1011_) );
      defparam ii1752.CONFIG_DATA = 16'h5555;
      defparam ii1752.PLACE_LOCATION = "NONE";
      defparam ii1752.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1753 ( .DX(nn1753), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1012_), .F2(dummy_abc_1013_), .F3(dummy_abc_1014_) );
      defparam ii1753.CONFIG_DATA = 16'h5555;
      defparam ii1753.PLACE_LOCATION = "NONE";
      defparam ii1753.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1754 ( .DX(nn1754), .F0(dummy_abc_1015_), .F1(dummy_abc_1016_), .F2(dummy_abc_1017_), .F3(dummy_abc_1018_) );
      defparam ii1754.CONFIG_DATA = 16'hFFFF;
      defparam ii1754.PLACE_LOCATION = "NONE";
      defparam ii1754.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_61_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_640_ ), 
        .DX( {nn1754, nn1753, nn1752, nn1751, nn1750, nn1749, nn1748, nn1747, 
              nn1746, nn1745, nn1744, nn1743, nn1742, nn1740, nn1738, nn1736, 
              nn1734, nn1733} ), 
        .SUM( {\coefcal1_divide_inst2_u130_XORCI_17|SUM_net , dummy_641_, 
              dummy_642_, dummy_643_, dummy_644_, dummy_645_, dummy_646_, dummy_647_, 
              dummy_648_, dummy_649_, dummy_650_, dummy_651_, dummy_652_, dummy_653_, 
              dummy_654_, dummy_655_, dummy_656_, dummy_657_} )
      );
    CS_LUT4_PRIM ii1775 ( .DX(nn1775), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1019_), .F3(dummy_abc_1020_) );
      defparam ii1775.CONFIG_DATA = 16'h9999;
      defparam ii1775.PLACE_LOCATION = "NONE";
      defparam ii1775.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1776 ( .DX(nn1776), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_640_) );
      defparam ii1776.CONFIG_DATA = 16'hA569;
      defparam ii1776.PLACE_LOCATION = "NONE";
      defparam ii1776.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1777 ( .DX(nn1777), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_621_), .F3(dummy_abc_1021_) );
      defparam ii1777.CONFIG_DATA = 16'hA6A6;
      defparam ii1777.PLACE_LOCATION = "NONE";
      defparam ii1777.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1778 ( .DX(nn1778), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1022_), .F3(dummy_abc_1023_) );
      defparam ii1778.CONFIG_DATA = 16'h9999;
      defparam ii1778.PLACE_LOCATION = "NONE";
      defparam ii1778.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1779 ( .DX(nn1779), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_621_) );
      defparam ii1779.CONFIG_DATA = 16'hA569;
      defparam ii1779.PLACE_LOCATION = "NONE";
      defparam ii1779.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1780 ( .DX(nn1780), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1735), .F2(dummy_abc_1024_), .F3(dummy_abc_1025_) );
      defparam ii1780.CONFIG_DATA = 16'h9999;
      defparam ii1780.PLACE_LOCATION = "NONE";
      defparam ii1780.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1781 ( .DX(nn1781), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1737), .F2(dummy_abc_1026_), .F3(dummy_abc_1027_) );
      defparam ii1781.CONFIG_DATA = 16'h9999;
      defparam ii1781.PLACE_LOCATION = "NONE";
      defparam ii1781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1782 ( .DX(nn1782), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1739), .F2(dummy_abc_1028_), .F3(dummy_abc_1029_) );
      defparam ii1782.CONFIG_DATA = 16'h9999;
      defparam ii1782.PLACE_LOCATION = "NONE";
      defparam ii1782.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1783 ( .DX(nn1783), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1741), .F2(dummy_abc_1030_), .F3(dummy_abc_1031_) );
      defparam ii1783.CONFIG_DATA = 16'h9999;
      defparam ii1783.PLACE_LOCATION = "NONE";
      defparam ii1783.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1784 ( .DX(nn1784), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1732), .F2(dummy_abc_1032_), .F3(dummy_abc_1033_) );
      defparam ii1784.CONFIG_DATA = 16'h9999;
      defparam ii1784.PLACE_LOCATION = "NONE";
      defparam ii1784.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1785 ( .DX(nn1785), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_1034_), .F2(dummy_abc_1035_), .F3(dummy_abc_1036_) );
      defparam ii1785.CONFIG_DATA = 16'h5555;
      defparam ii1785.PLACE_LOCATION = "NONE";
      defparam ii1785.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1786 ( .DX(nn1786), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1037_), .F2(dummy_abc_1038_), .F3(dummy_abc_1039_) );
      defparam ii1786.CONFIG_DATA = 16'h5555;
      defparam ii1786.PLACE_LOCATION = "NONE";
      defparam ii1786.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1787 ( .DX(nn1787), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1040_), .F2(dummy_abc_1041_), .F3(dummy_abc_1042_) );
      defparam ii1787.CONFIG_DATA = 16'h5555;
      defparam ii1787.PLACE_LOCATION = "NONE";
      defparam ii1787.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1788 ( .DX(nn1788), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1043_), .F2(dummy_abc_1044_), .F3(dummy_abc_1045_) );
      defparam ii1788.CONFIG_DATA = 16'h5555;
      defparam ii1788.PLACE_LOCATION = "NONE";
      defparam ii1788.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1789 ( .DX(nn1789), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1046_), .F2(dummy_abc_1047_), .F3(dummy_abc_1048_) );
      defparam ii1789.CONFIG_DATA = 16'h5555;
      defparam ii1789.PLACE_LOCATION = "NONE";
      defparam ii1789.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1790 ( .DX(nn1790), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1049_), .F2(dummy_abc_1050_), .F3(dummy_abc_1051_) );
      defparam ii1790.CONFIG_DATA = 16'h5555;
      defparam ii1790.PLACE_LOCATION = "NONE";
      defparam ii1790.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1791 ( .DX(nn1791), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1052_), .F2(dummy_abc_1053_), .F3(dummy_abc_1054_) );
      defparam ii1791.CONFIG_DATA = 16'h5555;
      defparam ii1791.PLACE_LOCATION = "NONE";
      defparam ii1791.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1792 ( .DX(nn1792), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1055_), .F2(dummy_abc_1056_), .F3(dummy_abc_1057_) );
      defparam ii1792.CONFIG_DATA = 16'h5555;
      defparam ii1792.PLACE_LOCATION = "NONE";
      defparam ii1792.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1793 ( .DX(nn1793), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1058_), .F2(dummy_abc_1059_), .F3(dummy_abc_1060_) );
      defparam ii1793.CONFIG_DATA = 16'h5555;
      defparam ii1793.PLACE_LOCATION = "NONE";
      defparam ii1793.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1794 ( .DX(nn1794), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1061_), .F2(dummy_abc_1062_), .F3(dummy_abc_1063_) );
      defparam ii1794.CONFIG_DATA = 16'h5555;
      defparam ii1794.PLACE_LOCATION = "NONE";
      defparam ii1794.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_45_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1732, nn1741, nn1739, nn1737, 
              nn1735, nn1777, \coefcal1_yDividend__reg[10]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_178_ ), 
        .DX( {nn1794, nn1793, nn1792, nn1791, nn1790, nn1789, nn1788, nn1787, 
              nn1786, nn1785, nn1784, nn1783, nn1782, nn1781, nn1780, nn1779, 
              nn1778} ), 
        .SUM( {dummy_179_, \coefcal1_divide_inst2_u107_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_14|SUM_net , \coefcal1_divide_inst2_u107_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_12|SUM_net , \coefcal1_divide_inst2_u107_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_10|SUM_net , \coefcal1_divide_inst2_u107_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_8|SUM_net , \coefcal1_divide_inst2_u107_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_6|SUM_net , \coefcal1_divide_inst2_u107_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_4|SUM_net , \coefcal1_divide_inst2_u107_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_2|SUM_net , \coefcal1_divide_inst2_u107_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1814 ( .DX(nn1814), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_640_), .F2(nn1777), .F3(\coefcal1_divide_inst2_u107_XORCI_1|SUM_net ) );
      defparam ii1814.CONFIG_DATA = 16'hA695;
      defparam ii1814.PLACE_LOCATION = "NONE";
      defparam ii1814.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1815 ( .DX(nn1815), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1735), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_2|SUM_net ) );
      defparam ii1815.CONFIG_DATA = 16'h9A95;
      defparam ii1815.PLACE_LOCATION = "NONE";
      defparam ii1815.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1816 ( .DX(nn1816), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1737), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_3|SUM_net ) );
      defparam ii1816.CONFIG_DATA = 16'h9A95;
      defparam ii1816.PLACE_LOCATION = "NONE";
      defparam ii1816.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1817 ( .DX(nn1817), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1739), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_4|SUM_net ) );
      defparam ii1817.CONFIG_DATA = 16'h9A95;
      defparam ii1817.PLACE_LOCATION = "NONE";
      defparam ii1817.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1818 ( .DX(nn1818), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1741), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_5|SUM_net ) );
      defparam ii1818.CONFIG_DATA = 16'h9A95;
      defparam ii1818.PLACE_LOCATION = "NONE";
      defparam ii1818.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1819 ( .DX(nn1819), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1732), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_6|SUM_net ) );
      defparam ii1819.CONFIG_DATA = 16'h9A95;
      defparam ii1819.PLACE_LOCATION = "NONE";
      defparam ii1819.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1820 ( .DX(nn1820), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1064_), .F2(dummy_abc_1065_), .F3(dummy_abc_1066_) );
      defparam ii1820.CONFIG_DATA = 16'h5555;
      defparam ii1820.PLACE_LOCATION = "NONE";
      defparam ii1820.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1821 ( .DX(nn1821), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1067_), .F2(dummy_abc_1068_), .F3(dummy_abc_1069_) );
      defparam ii1821.CONFIG_DATA = 16'h5555;
      defparam ii1821.PLACE_LOCATION = "NONE";
      defparam ii1821.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1822 ( .DX(nn1822), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1070_), .F2(dummy_abc_1071_), .F3(dummy_abc_1072_) );
      defparam ii1822.CONFIG_DATA = 16'h5555;
      defparam ii1822.PLACE_LOCATION = "NONE";
      defparam ii1822.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1823 ( .DX(nn1823), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1073_), .F2(dummy_abc_1074_), .F3(dummy_abc_1075_) );
      defparam ii1823.CONFIG_DATA = 16'h5555;
      defparam ii1823.PLACE_LOCATION = "NONE";
      defparam ii1823.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1824 ( .DX(nn1824), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1076_), .F2(dummy_abc_1077_), .F3(dummy_abc_1078_) );
      defparam ii1824.CONFIG_DATA = 16'h5555;
      defparam ii1824.PLACE_LOCATION = "NONE";
      defparam ii1824.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1825 ( .DX(nn1825), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1079_), .F2(dummy_abc_1080_), .F3(dummy_abc_1081_) );
      defparam ii1825.CONFIG_DATA = 16'h5555;
      defparam ii1825.PLACE_LOCATION = "NONE";
      defparam ii1825.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1826 ( .DX(nn1826), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1082_), .F2(dummy_abc_1083_), .F3(dummy_abc_1084_) );
      defparam ii1826.CONFIG_DATA = 16'h5555;
      defparam ii1826.PLACE_LOCATION = "NONE";
      defparam ii1826.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1827 ( .DX(nn1827), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1085_), .F2(dummy_abc_1086_), .F3(dummy_abc_1087_) );
      defparam ii1827.CONFIG_DATA = 16'h5555;
      defparam ii1827.PLACE_LOCATION = "NONE";
      defparam ii1827.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1828 ( .DX(nn1828), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1088_), .F2(dummy_abc_1089_), .F3(dummy_abc_1090_) );
      defparam ii1828.CONFIG_DATA = 16'h5555;
      defparam ii1828.PLACE_LOCATION = "NONE";
      defparam ii1828.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1829 ( .DX(nn1829), .F0(dummy_abc_1091_), .F1(dummy_abc_1092_), .F2(dummy_abc_1093_), .F3(dummy_abc_1094_) );
      defparam ii1829.CONFIG_DATA = 16'hFFFF;
      defparam ii1829.PLACE_LOCATION = "NONE";
      defparam ii1829.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_62_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_659_ ), 
        .DX( {nn1829, nn1828, nn1827, nn1826, nn1825, nn1824, nn1823, nn1822, 
              nn1821, nn1820, nn1819, nn1818, nn1817, nn1816, nn1815, nn1814, 
              nn1776, nn1775} ), 
        .SUM( {\coefcal1_divide_inst2_u132_XORCI_17|SUM_net , dummy_660_, 
              dummy_661_, dummy_662_, dummy_663_, dummy_664_, dummy_665_, dummy_666_, 
              dummy_667_, dummy_668_, dummy_669_, dummy_670_, dummy_671_, dummy_672_, 
              dummy_673_, dummy_674_, dummy_675_, dummy_676_} )
      );
    CS_LUT4_PRIM ii1850 ( .DX(nn1850), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_640_), .F3(dummy_abc_1095_) );
      defparam ii1850.CONFIG_DATA = 16'hA6A6;
      defparam ii1850.PLACE_LOCATION = "NONE";
      defparam ii1850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1851 ( .DX(nn1851), .F0(dummy_640_), .F1(nn1777), .F2(\coefcal1_divide_inst2_u107_XORCI_1|SUM_net ), .F3(dummy_abc_1096_) );
      defparam ii1851.CONFIG_DATA = 16'hD8D8;
      defparam ii1851.PLACE_LOCATION = "NONE";
      defparam ii1851.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1852 ( .DX(nn1852), .F0(nn1735), .F1(dummy_640_), .F2(\coefcal1_divide_inst2_u107_XORCI_2|SUM_net ), .F3(dummy_abc_1097_) );
      defparam ii1852.CONFIG_DATA = 16'hB8B8;
      defparam ii1852.PLACE_LOCATION = "NONE";
      defparam ii1852.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1853 ( .DX(nn1853), .F0(nn1737), .F1(dummy_640_), .F2(\coefcal1_divide_inst2_u107_XORCI_3|SUM_net ), .F3(dummy_abc_1098_) );
      defparam ii1853.CONFIG_DATA = 16'hB8B8;
      defparam ii1853.PLACE_LOCATION = "NONE";
      defparam ii1853.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1854 ( .DX(nn1854), .F0(nn1739), .F1(dummy_640_), .F2(\coefcal1_divide_inst2_u107_XORCI_4|SUM_net ), .F3(dummy_abc_1099_) );
      defparam ii1854.CONFIG_DATA = 16'hB8B8;
      defparam ii1854.PLACE_LOCATION = "NONE";
      defparam ii1854.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1855 ( .DX(nn1855), .F0(nn1741), .F1(dummy_640_), .F2(\coefcal1_divide_inst2_u107_XORCI_5|SUM_net ), .F3(dummy_abc_1100_) );
      defparam ii1855.CONFIG_DATA = 16'hB8B8;
      defparam ii1855.PLACE_LOCATION = "NONE";
      defparam ii1855.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1856 ( .DX(nn1856), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1101_), .F3(dummy_abc_1102_) );
      defparam ii1856.CONFIG_DATA = 16'h9999;
      defparam ii1856.PLACE_LOCATION = "NONE";
      defparam ii1856.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1857 ( .DX(nn1857), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_640_) );
      defparam ii1857.CONFIG_DATA = 16'hA569;
      defparam ii1857.PLACE_LOCATION = "NONE";
      defparam ii1857.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1858 ( .DX(nn1858), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_640_), .F2(nn1777), .F3(\coefcal1_divide_inst2_u107_XORCI_1|SUM_net ) );
      defparam ii1858.CONFIG_DATA = 16'hA695;
      defparam ii1858.PLACE_LOCATION = "NONE";
      defparam ii1858.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1859 ( .DX(nn1859), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1735), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_2|SUM_net ) );
      defparam ii1859.CONFIG_DATA = 16'h9A95;
      defparam ii1859.PLACE_LOCATION = "NONE";
      defparam ii1859.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1860 ( .DX(nn1860), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1737), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_3|SUM_net ) );
      defparam ii1860.CONFIG_DATA = 16'h9A95;
      defparam ii1860.PLACE_LOCATION = "NONE";
      defparam ii1860.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1861 ( .DX(nn1861), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1739), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_4|SUM_net ) );
      defparam ii1861.CONFIG_DATA = 16'h9A95;
      defparam ii1861.PLACE_LOCATION = "NONE";
      defparam ii1861.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1862 ( .DX(nn1862), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1741), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_5|SUM_net ) );
      defparam ii1862.CONFIG_DATA = 16'h9A95;
      defparam ii1862.PLACE_LOCATION = "NONE";
      defparam ii1862.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1863 ( .DX(nn1863), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1732), .F2(dummy_640_), .F3(\coefcal1_divide_inst2_u107_XORCI_6|SUM_net ) );
      defparam ii1863.CONFIG_DATA = 16'h9A95;
      defparam ii1863.PLACE_LOCATION = "NONE";
      defparam ii1863.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1864 ( .DX(nn1864), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1103_), .F2(dummy_abc_1104_), .F3(dummy_abc_1105_) );
      defparam ii1864.CONFIG_DATA = 16'h5555;
      defparam ii1864.PLACE_LOCATION = "NONE";
      defparam ii1864.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1865 ( .DX(nn1865), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1106_), .F2(dummy_abc_1107_), .F3(dummy_abc_1108_) );
      defparam ii1865.CONFIG_DATA = 16'h5555;
      defparam ii1865.PLACE_LOCATION = "NONE";
      defparam ii1865.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1866 ( .DX(nn1866), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1109_), .F2(dummy_abc_1110_), .F3(dummy_abc_1111_) );
      defparam ii1866.CONFIG_DATA = 16'h5555;
      defparam ii1866.PLACE_LOCATION = "NONE";
      defparam ii1866.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1867 ( .DX(nn1867), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1112_), .F2(dummy_abc_1113_), .F3(dummy_abc_1114_) );
      defparam ii1867.CONFIG_DATA = 16'h5555;
      defparam ii1867.PLACE_LOCATION = "NONE";
      defparam ii1867.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1868 ( .DX(nn1868), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1115_), .F2(dummy_abc_1116_), .F3(dummy_abc_1117_) );
      defparam ii1868.CONFIG_DATA = 16'h5555;
      defparam ii1868.PLACE_LOCATION = "NONE";
      defparam ii1868.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1869 ( .DX(nn1869), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1118_), .F2(dummy_abc_1119_), .F3(dummy_abc_1120_) );
      defparam ii1869.CONFIG_DATA = 16'h5555;
      defparam ii1869.PLACE_LOCATION = "NONE";
      defparam ii1869.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1870 ( .DX(nn1870), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1121_), .F2(dummy_abc_1122_), .F3(dummy_abc_1123_) );
      defparam ii1870.CONFIG_DATA = 16'h5555;
      defparam ii1870.PLACE_LOCATION = "NONE";
      defparam ii1870.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1871 ( .DX(nn1871), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1124_), .F2(dummy_abc_1125_), .F3(dummy_abc_1126_) );
      defparam ii1871.CONFIG_DATA = 16'h5555;
      defparam ii1871.PLACE_LOCATION = "NONE";
      defparam ii1871.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1872 ( .DX(nn1872), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1127_), .F2(dummy_abc_1128_), .F3(dummy_abc_1129_) );
      defparam ii1872.CONFIG_DATA = 16'h5555;
      defparam ii1872.PLACE_LOCATION = "NONE";
      defparam ii1872.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_46_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1855, nn1854, nn1853, nn1852, 
              nn1851, nn1850, \coefcal1_yDividend__reg[9]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_180_ ), 
        .DX( {nn1872, nn1871, nn1870, nn1869, nn1868, nn1867, nn1866, nn1865, 
              nn1864, nn1863, nn1862, nn1861, nn1860, nn1859, nn1858, nn1857, 
              nn1856} ), 
        .SUM( {dummy_181_, \coefcal1_divide_inst2_u108_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_14|SUM_net , \coefcal1_divide_inst2_u108_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_12|SUM_net , \coefcal1_divide_inst2_u108_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_10|SUM_net , \coefcal1_divide_inst2_u108_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_8|SUM_net , \coefcal1_divide_inst2_u108_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_6|SUM_net , \coefcal1_divide_inst2_u108_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_4|SUM_net , \coefcal1_divide_inst2_u108_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_2|SUM_net , \coefcal1_divide_inst2_u108_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1892 ( .DX(nn1892), .F0(nn1732), .F1(dummy_640_), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ) );
      defparam ii1892.CONFIG_DATA = 16'h8F80;
      defparam ii1892.PLACE_LOCATION = "NONE";
      defparam ii1892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1893 ( .DX(nn1893), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1130_), .F3(dummy_abc_1131_) );
      defparam ii1893.CONFIG_DATA = 16'h9999;
      defparam ii1893.PLACE_LOCATION = "NONE";
      defparam ii1893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1894 ( .DX(nn1894), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_659_) );
      defparam ii1894.CONFIG_DATA = 16'hA569;
      defparam ii1894.PLACE_LOCATION = "NONE";
      defparam ii1894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1895 ( .DX(nn1895), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_659_), .F2(nn1850), .F3(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ) );
      defparam ii1895.CONFIG_DATA = 16'hA695;
      defparam ii1895.PLACE_LOCATION = "NONE";
      defparam ii1895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1896 ( .DX(nn1896), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1851), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ) );
      defparam ii1896.CONFIG_DATA = 16'h9A95;
      defparam ii1896.PLACE_LOCATION = "NONE";
      defparam ii1896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1897 ( .DX(nn1897), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1852), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ) );
      defparam ii1897.CONFIG_DATA = 16'h9A95;
      defparam ii1897.PLACE_LOCATION = "NONE";
      defparam ii1897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1898 ( .DX(nn1898), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1853), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ) );
      defparam ii1898.CONFIG_DATA = 16'h9A95;
      defparam ii1898.PLACE_LOCATION = "NONE";
      defparam ii1898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1899 ( .DX(nn1899), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1854), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ) );
      defparam ii1899.CONFIG_DATA = 16'h9A95;
      defparam ii1899.PLACE_LOCATION = "NONE";
      defparam ii1899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1900 ( .DX(nn1900), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1855), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ) );
      defparam ii1900.CONFIG_DATA = 16'h9A95;
      defparam ii1900.PLACE_LOCATION = "NONE";
      defparam ii1900.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1901 ( .DX(nn1901), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn1732), .F2(dummy_640_), .F3(dummy_abc_1132_) );
      defparam ii1901.CONFIG_DATA = 16'h9595;
      defparam ii1901.PLACE_LOCATION = "NONE";
      defparam ii1901.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1902 ( .DX(nn1902), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ), .F3(nn1901) );
      defparam ii1902.CONFIG_DATA = 16'hCD01;
      defparam ii1902.PLACE_LOCATION = "NONE";
      defparam ii1902.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1903 ( .DX(nn1903), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1133_), .F2(dummy_abc_1134_), .F3(dummy_abc_1135_) );
      defparam ii1903.CONFIG_DATA = 16'h5555;
      defparam ii1903.PLACE_LOCATION = "NONE";
      defparam ii1903.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1904 ( .DX(nn1904), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1136_), .F2(dummy_abc_1137_), .F3(dummy_abc_1138_) );
      defparam ii1904.CONFIG_DATA = 16'h5555;
      defparam ii1904.PLACE_LOCATION = "NONE";
      defparam ii1904.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1905 ( .DX(nn1905), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1139_), .F2(dummy_abc_1140_), .F3(dummy_abc_1141_) );
      defparam ii1905.CONFIG_DATA = 16'h5555;
      defparam ii1905.PLACE_LOCATION = "NONE";
      defparam ii1905.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1906 ( .DX(nn1906), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1142_), .F2(dummy_abc_1143_), .F3(dummy_abc_1144_) );
      defparam ii1906.CONFIG_DATA = 16'h5555;
      defparam ii1906.PLACE_LOCATION = "NONE";
      defparam ii1906.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1907 ( .DX(nn1907), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1145_), .F2(dummy_abc_1146_), .F3(dummy_abc_1147_) );
      defparam ii1907.CONFIG_DATA = 16'h5555;
      defparam ii1907.PLACE_LOCATION = "NONE";
      defparam ii1907.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1908 ( .DX(nn1908), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1148_), .F2(dummy_abc_1149_), .F3(dummy_abc_1150_) );
      defparam ii1908.CONFIG_DATA = 16'h5555;
      defparam ii1908.PLACE_LOCATION = "NONE";
      defparam ii1908.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1909 ( .DX(nn1909), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1151_), .F2(dummy_abc_1152_), .F3(dummy_abc_1153_) );
      defparam ii1909.CONFIG_DATA = 16'h5555;
      defparam ii1909.PLACE_LOCATION = "NONE";
      defparam ii1909.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1910 ( .DX(nn1910), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1154_), .F2(dummy_abc_1155_), .F3(dummy_abc_1156_) );
      defparam ii1910.CONFIG_DATA = 16'h5555;
      defparam ii1910.PLACE_LOCATION = "NONE";
      defparam ii1910.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1911 ( .DX(nn1911), .F0(dummy_abc_1157_), .F1(dummy_abc_1158_), .F2(dummy_abc_1159_), .F3(dummy_abc_1160_) );
      defparam ii1911.CONFIG_DATA = 16'hFFFF;
      defparam ii1911.PLACE_LOCATION = "NONE";
      defparam ii1911.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_63_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_678_ ), 
        .DX( {nn1911, nn1910, nn1909, nn1908, nn1907, nn1906, nn1905, nn1904, 
              nn1903, nn1902, nn1900, nn1899, nn1898, nn1897, nn1896, nn1895, 
              nn1894, nn1893} ), 
        .SUM( {\coefcal1_divide_inst2_u134_XORCI_17|SUM_net , dummy_679_, 
              dummy_680_, dummy_681_, dummy_682_, dummy_683_, dummy_684_, dummy_685_, 
              dummy_686_, dummy_687_, dummy_688_, dummy_689_, dummy_690_, dummy_691_, 
              dummy_692_, dummy_693_, dummy_694_, dummy_695_} )
      );
    CS_LUT4_PRIM ii1932 ( .DX(nn1932), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_659_), .F3(dummy_abc_1161_) );
      defparam ii1932.CONFIG_DATA = 16'hA6A6;
      defparam ii1932.PLACE_LOCATION = "NONE";
      defparam ii1932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1933 ( .DX(nn1933), .F0(dummy_659_), .F1(nn1850), .F2(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ), .F3(dummy_abc_1162_) );
      defparam ii1933.CONFIG_DATA = 16'hD8D8;
      defparam ii1933.PLACE_LOCATION = "NONE";
      defparam ii1933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1934 ( .DX(nn1934), .F0(nn1851), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ), .F3(dummy_abc_1163_) );
      defparam ii1934.CONFIG_DATA = 16'hB8B8;
      defparam ii1934.PLACE_LOCATION = "NONE";
      defparam ii1934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1935 ( .DX(nn1935), .F0(nn1852), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ), .F3(dummy_abc_1164_) );
      defparam ii1935.CONFIG_DATA = 16'hB8B8;
      defparam ii1935.PLACE_LOCATION = "NONE";
      defparam ii1935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1936 ( .DX(nn1936), .F0(nn1853), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ), .F3(dummy_abc_1165_) );
      defparam ii1936.CONFIG_DATA = 16'hB8B8;
      defparam ii1936.PLACE_LOCATION = "NONE";
      defparam ii1936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1937 ( .DX(nn1937), .F0(nn1854), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ), .F3(dummy_abc_1166_) );
      defparam ii1937.CONFIG_DATA = 16'hB8B8;
      defparam ii1937.PLACE_LOCATION = "NONE";
      defparam ii1937.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1938 ( .DX(nn1938), .F0(nn1855), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ), .F3(dummy_abc_1167_) );
      defparam ii1938.CONFIG_DATA = 16'hB8B8;
      defparam ii1938.PLACE_LOCATION = "NONE";
      defparam ii1938.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1939 ( .DX(nn1939), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1168_), .F3(dummy_abc_1169_) );
      defparam ii1939.CONFIG_DATA = 16'h9999;
      defparam ii1939.PLACE_LOCATION = "NONE";
      defparam ii1939.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1940 ( .DX(nn1940), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_659_) );
      defparam ii1940.CONFIG_DATA = 16'hA569;
      defparam ii1940.PLACE_LOCATION = "NONE";
      defparam ii1940.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1941 ( .DX(nn1941), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_659_), .F2(nn1850), .F3(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ) );
      defparam ii1941.CONFIG_DATA = 16'hA695;
      defparam ii1941.PLACE_LOCATION = "NONE";
      defparam ii1941.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1942 ( .DX(nn1942), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1851), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ) );
      defparam ii1942.CONFIG_DATA = 16'h9A95;
      defparam ii1942.PLACE_LOCATION = "NONE";
      defparam ii1942.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1943 ( .DX(nn1943), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1852), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ) );
      defparam ii1943.CONFIG_DATA = 16'h9A95;
      defparam ii1943.PLACE_LOCATION = "NONE";
      defparam ii1943.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1944 ( .DX(nn1944), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1853), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ) );
      defparam ii1944.CONFIG_DATA = 16'h9A95;
      defparam ii1944.PLACE_LOCATION = "NONE";
      defparam ii1944.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1945 ( .DX(nn1945), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1854), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ) );
      defparam ii1945.CONFIG_DATA = 16'h9A95;
      defparam ii1945.PLACE_LOCATION = "NONE";
      defparam ii1945.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1946 ( .DX(nn1946), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1855), .F2(dummy_659_), .F3(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ) );
      defparam ii1946.CONFIG_DATA = 16'h9A95;
      defparam ii1946.PLACE_LOCATION = "NONE";
      defparam ii1946.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1947 ( .DX(nn1947), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_659_), .F2(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ), .F3(nn1901) );
      defparam ii1947.CONFIG_DATA = 16'hCD01;
      defparam ii1947.PLACE_LOCATION = "NONE";
      defparam ii1947.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1948 ( .DX(nn1948), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1170_), .F2(dummy_abc_1171_), .F3(dummy_abc_1172_) );
      defparam ii1948.CONFIG_DATA = 16'h5555;
      defparam ii1948.PLACE_LOCATION = "NONE";
      defparam ii1948.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1949 ( .DX(nn1949), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1173_), .F2(dummy_abc_1174_), .F3(dummy_abc_1175_) );
      defparam ii1949.CONFIG_DATA = 16'h5555;
      defparam ii1949.PLACE_LOCATION = "NONE";
      defparam ii1949.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1950 ( .DX(nn1950), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1176_), .F2(dummy_abc_1177_), .F3(dummy_abc_1178_) );
      defparam ii1950.CONFIG_DATA = 16'h5555;
      defparam ii1950.PLACE_LOCATION = "NONE";
      defparam ii1950.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1951 ( .DX(nn1951), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1179_), .F2(dummy_abc_1180_), .F3(dummy_abc_1181_) );
      defparam ii1951.CONFIG_DATA = 16'h5555;
      defparam ii1951.PLACE_LOCATION = "NONE";
      defparam ii1951.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1952 ( .DX(nn1952), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1182_), .F2(dummy_abc_1183_), .F3(dummy_abc_1184_) );
      defparam ii1952.CONFIG_DATA = 16'h5555;
      defparam ii1952.PLACE_LOCATION = "NONE";
      defparam ii1952.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1953 ( .DX(nn1953), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1185_), .F2(dummy_abc_1186_), .F3(dummy_abc_1187_) );
      defparam ii1953.CONFIG_DATA = 16'h5555;
      defparam ii1953.PLACE_LOCATION = "NONE";
      defparam ii1953.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1954 ( .DX(nn1954), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1188_), .F2(dummy_abc_1189_), .F3(dummy_abc_1190_) );
      defparam ii1954.CONFIG_DATA = 16'h5555;
      defparam ii1954.PLACE_LOCATION = "NONE";
      defparam ii1954.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1955 ( .DX(nn1955), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1191_), .F2(dummy_abc_1192_), .F3(dummy_abc_1193_) );
      defparam ii1955.CONFIG_DATA = 16'h5555;
      defparam ii1955.PLACE_LOCATION = "NONE";
      defparam ii1955.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_47_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn1892, 
              nn1938, nn1937, nn1936, nn1935, nn1934, nn1933, nn1932, 
              \coefcal1_yDividend__reg[8]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_182_ ), 
        .DX( {nn1955, nn1954, nn1953, nn1952, nn1951, nn1950, nn1949, nn1948, 
              nn1947, nn1946, nn1945, nn1944, nn1943, nn1942, nn1941, nn1940, 
              nn1939} ), 
        .SUM( {dummy_183_, \coefcal1_divide_inst2_u109_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_14|SUM_net , \coefcal1_divide_inst2_u109_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_12|SUM_net , \coefcal1_divide_inst2_u109_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_10|SUM_net , \coefcal1_divide_inst2_u109_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_8|SUM_net , \coefcal1_divide_inst2_u109_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_6|SUM_net , \coefcal1_divide_inst2_u109_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_4|SUM_net , \coefcal1_divide_inst2_u109_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_2|SUM_net , \coefcal1_divide_inst2_u109_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1975 ( .DX(nn1975), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1194_), .F3(dummy_abc_1195_) );
      defparam ii1975.CONFIG_DATA = 16'h9999;
      defparam ii1975.PLACE_LOCATION = "NONE";
      defparam ii1975.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1976 ( .DX(nn1976), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_678_) );
      defparam ii1976.CONFIG_DATA = 16'hA569;
      defparam ii1976.PLACE_LOCATION = "NONE";
      defparam ii1976.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1977 ( .DX(nn1977), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_678_), .F2(nn1932), .F3(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ) );
      defparam ii1977.CONFIG_DATA = 16'hA695;
      defparam ii1977.PLACE_LOCATION = "NONE";
      defparam ii1977.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1978 ( .DX(nn1978), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1933), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ) );
      defparam ii1978.CONFIG_DATA = 16'h9A95;
      defparam ii1978.PLACE_LOCATION = "NONE";
      defparam ii1978.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1979 ( .DX(nn1979), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1934), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ) );
      defparam ii1979.CONFIG_DATA = 16'h9A95;
      defparam ii1979.PLACE_LOCATION = "NONE";
      defparam ii1979.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1980 ( .DX(nn1980), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1935), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ) );
      defparam ii1980.CONFIG_DATA = 16'h9A95;
      defparam ii1980.PLACE_LOCATION = "NONE";
      defparam ii1980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1981 ( .DX(nn1981), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1936), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ) );
      defparam ii1981.CONFIG_DATA = 16'h9A95;
      defparam ii1981.PLACE_LOCATION = "NONE";
      defparam ii1981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1982 ( .DX(nn1982), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1937), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ) );
      defparam ii1982.CONFIG_DATA = 16'h9A95;
      defparam ii1982.PLACE_LOCATION = "NONE";
      defparam ii1982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1983 ( .DX(nn1983), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn1938), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ) );
      defparam ii1983.CONFIG_DATA = 16'h9A95;
      defparam ii1983.PLACE_LOCATION = "NONE";
      defparam ii1983.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1984 ( .DX(nn1984), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn1892), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ) );
      defparam ii1984.CONFIG_DATA = 16'h9995;
      defparam ii1984.PLACE_LOCATION = "NONE";
      defparam ii1984.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1985 ( .DX(nn1985), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1196_), .F2(dummy_abc_1197_), .F3(dummy_abc_1198_) );
      defparam ii1985.CONFIG_DATA = 16'h5555;
      defparam ii1985.PLACE_LOCATION = "NONE";
      defparam ii1985.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1986 ( .DX(nn1986), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1199_), .F2(dummy_abc_1200_), .F3(dummy_abc_1201_) );
      defparam ii1986.CONFIG_DATA = 16'h5555;
      defparam ii1986.PLACE_LOCATION = "NONE";
      defparam ii1986.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1987 ( .DX(nn1987), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1202_), .F2(dummy_abc_1203_), .F3(dummy_abc_1204_) );
      defparam ii1987.CONFIG_DATA = 16'h5555;
      defparam ii1987.PLACE_LOCATION = "NONE";
      defparam ii1987.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1988 ( .DX(nn1988), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1205_), .F2(dummy_abc_1206_), .F3(dummy_abc_1207_) );
      defparam ii1988.CONFIG_DATA = 16'h5555;
      defparam ii1988.PLACE_LOCATION = "NONE";
      defparam ii1988.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1989 ( .DX(nn1989), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1208_), .F2(dummy_abc_1209_), .F3(dummy_abc_1210_) );
      defparam ii1989.CONFIG_DATA = 16'h5555;
      defparam ii1989.PLACE_LOCATION = "NONE";
      defparam ii1989.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1990 ( .DX(nn1990), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1211_), .F2(dummy_abc_1212_), .F3(dummy_abc_1213_) );
      defparam ii1990.CONFIG_DATA = 16'h5555;
      defparam ii1990.PLACE_LOCATION = "NONE";
      defparam ii1990.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1991 ( .DX(nn1991), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1214_), .F2(dummy_abc_1215_), .F3(dummy_abc_1216_) );
      defparam ii1991.CONFIG_DATA = 16'h5555;
      defparam ii1991.PLACE_LOCATION = "NONE";
      defparam ii1991.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1992 ( .DX(nn1992), .F0(dummy_abc_1217_), .F1(dummy_abc_1218_), .F2(dummy_abc_1219_), .F3(dummy_abc_1220_) );
      defparam ii1992.CONFIG_DATA = 16'hFFFF;
      defparam ii1992.PLACE_LOCATION = "NONE";
      defparam ii1992.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_64_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_697_ ), 
        .DX( {nn1992, nn1991, nn1990, nn1989, nn1988, nn1987, nn1986, nn1985, 
              nn1984, nn1983, nn1982, nn1981, nn1980, nn1979, nn1978, nn1977, 
              nn1976, nn1975} ), 
        .SUM( {\coefcal1_divide_inst2_u136_XORCI_17|SUM_net , dummy_698_, 
              dummy_699_, dummy_700_, dummy_701_, dummy_702_, dummy_703_, dummy_704_, 
              dummy_705_, dummy_706_, dummy_707_, dummy_708_, dummy_709_, dummy_710_, 
              dummy_711_, dummy_712_, dummy_713_, dummy_714_} )
      );
    CS_LUT4_PRIM ii2013 ( .DX(nn2013), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_678_), .F3(dummy_abc_1221_) );
      defparam ii2013.CONFIG_DATA = 16'hA6A6;
      defparam ii2013.PLACE_LOCATION = "NONE";
      defparam ii2013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2014 ( .DX(nn2014), .F0(dummy_678_), .F1(nn1932), .F2(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ), .F3(dummy_abc_1222_) );
      defparam ii2014.CONFIG_DATA = 16'hD8D8;
      defparam ii2014.PLACE_LOCATION = "NONE";
      defparam ii2014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2015 ( .DX(nn2015), .F0(nn1933), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ), .F3(dummy_abc_1223_) );
      defparam ii2015.CONFIG_DATA = 16'hB8B8;
      defparam ii2015.PLACE_LOCATION = "NONE";
      defparam ii2015.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2016 ( .DX(nn2016), .F0(nn1934), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ), .F3(dummy_abc_1224_) );
      defparam ii2016.CONFIG_DATA = 16'hB8B8;
      defparam ii2016.PLACE_LOCATION = "NONE";
      defparam ii2016.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2017 ( .DX(nn2017), .F0(nn1935), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ), .F3(dummy_abc_1225_) );
      defparam ii2017.CONFIG_DATA = 16'hB8B8;
      defparam ii2017.PLACE_LOCATION = "NONE";
      defparam ii2017.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2018 ( .DX(nn2018), .F0(nn1936), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ), .F3(dummy_abc_1226_) );
      defparam ii2018.CONFIG_DATA = 16'hB8B8;
      defparam ii2018.PLACE_LOCATION = "NONE";
      defparam ii2018.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2019 ( .DX(nn2019), .F0(nn1937), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ), .F3(dummy_abc_1227_) );
      defparam ii2019.CONFIG_DATA = 16'hB8B8;
      defparam ii2019.PLACE_LOCATION = "NONE";
      defparam ii2019.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2020 ( .DX(nn2020), .F0(nn1938), .F1(dummy_678_), .F2(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ), .F3(dummy_abc_1228_) );
      defparam ii2020.CONFIG_DATA = 16'hB8B8;
      defparam ii2020.PLACE_LOCATION = "NONE";
      defparam ii2020.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2021 ( .DX(nn2021), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1229_), .F3(dummy_abc_1230_) );
      defparam ii2021.CONFIG_DATA = 16'h9999;
      defparam ii2021.PLACE_LOCATION = "NONE";
      defparam ii2021.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2022 ( .DX(nn2022), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_678_) );
      defparam ii2022.CONFIG_DATA = 16'hA569;
      defparam ii2022.PLACE_LOCATION = "NONE";
      defparam ii2022.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2023 ( .DX(nn2023), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_678_), .F2(nn1932), .F3(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ) );
      defparam ii2023.CONFIG_DATA = 16'hA695;
      defparam ii2023.PLACE_LOCATION = "NONE";
      defparam ii2023.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2024 ( .DX(nn2024), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1933), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ) );
      defparam ii2024.CONFIG_DATA = 16'h9A95;
      defparam ii2024.PLACE_LOCATION = "NONE";
      defparam ii2024.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2025 ( .DX(nn2025), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1934), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ) );
      defparam ii2025.CONFIG_DATA = 16'h9A95;
      defparam ii2025.PLACE_LOCATION = "NONE";
      defparam ii2025.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2026 ( .DX(nn2026), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1935), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ) );
      defparam ii2026.CONFIG_DATA = 16'h9A95;
      defparam ii2026.PLACE_LOCATION = "NONE";
      defparam ii2026.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2027 ( .DX(nn2027), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1936), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ) );
      defparam ii2027.CONFIG_DATA = 16'h9A95;
      defparam ii2027.PLACE_LOCATION = "NONE";
      defparam ii2027.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2028 ( .DX(nn2028), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1937), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ) );
      defparam ii2028.CONFIG_DATA = 16'h9A95;
      defparam ii2028.PLACE_LOCATION = "NONE";
      defparam ii2028.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2029 ( .DX(nn2029), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn1938), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ) );
      defparam ii2029.CONFIG_DATA = 16'h9A95;
      defparam ii2029.PLACE_LOCATION = "NONE";
      defparam ii2029.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2030 ( .DX(nn2030), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn1892), .F2(dummy_678_), .F3(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ) );
      defparam ii2030.CONFIG_DATA = 16'h9995;
      defparam ii2030.PLACE_LOCATION = "NONE";
      defparam ii2030.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2031 ( .DX(nn2031), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1231_), .F2(dummy_abc_1232_), .F3(dummy_abc_1233_) );
      defparam ii2031.CONFIG_DATA = 16'h5555;
      defparam ii2031.PLACE_LOCATION = "NONE";
      defparam ii2031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2032 ( .DX(nn2032), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1234_), .F2(dummy_abc_1235_), .F3(dummy_abc_1236_) );
      defparam ii2032.CONFIG_DATA = 16'h5555;
      defparam ii2032.PLACE_LOCATION = "NONE";
      defparam ii2032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2033 ( .DX(nn2033), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1237_), .F2(dummy_abc_1238_), .F3(dummy_abc_1239_) );
      defparam ii2033.CONFIG_DATA = 16'h5555;
      defparam ii2033.PLACE_LOCATION = "NONE";
      defparam ii2033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2034 ( .DX(nn2034), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1240_), .F2(dummy_abc_1241_), .F3(dummy_abc_1242_) );
      defparam ii2034.CONFIG_DATA = 16'h5555;
      defparam ii2034.PLACE_LOCATION = "NONE";
      defparam ii2034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2035 ( .DX(nn2035), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1243_), .F2(dummy_abc_1244_), .F3(dummy_abc_1245_) );
      defparam ii2035.CONFIG_DATA = 16'h5555;
      defparam ii2035.PLACE_LOCATION = "NONE";
      defparam ii2035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2036 ( .DX(nn2036), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1246_), .F2(dummy_abc_1247_), .F3(dummy_abc_1248_) );
      defparam ii2036.CONFIG_DATA = 16'h5555;
      defparam ii2036.PLACE_LOCATION = "NONE";
      defparam ii2036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2037 ( .DX(nn2037), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1249_), .F2(dummy_abc_1250_), .F3(dummy_abc_1251_) );
      defparam ii2037.CONFIG_DATA = 16'h5555;
      defparam ii2037.PLACE_LOCATION = "NONE";
      defparam ii2037.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_48_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2020, 
              nn2019, nn2018, nn2017, nn2016, nn2015, nn2014, nn2013, 
              \coefcal1_yDividend__reg[7]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_184_ ), 
        .DX( {nn2037, nn2036, nn2035, nn2034, nn2033, nn2032, nn2031, nn2030, 
              nn2029, nn2028, nn2027, nn2026, nn2025, nn2024, nn2023, nn2022, 
              nn2021} ), 
        .SUM( {dummy_185_, \coefcal1_divide_inst2_u110_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_14|SUM_net , \coefcal1_divide_inst2_u110_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_12|SUM_net , \coefcal1_divide_inst2_u110_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_10|SUM_net , \coefcal1_divide_inst2_u110_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_8|SUM_net , \coefcal1_divide_inst2_u110_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_6|SUM_net , \coefcal1_divide_inst2_u110_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_4|SUM_net , \coefcal1_divide_inst2_u110_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_2|SUM_net , \coefcal1_divide_inst2_u110_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2057 ( .DX(nn2057), .F0(dummy_678_), .F1(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ), .F2(dummy_697_), .F3(\coefcal1_divide_inst2_u110_XORCI_9|SUM_net ) );
      defparam ii2057.CONFIG_DATA = 16'hEFE0;
      defparam ii2057.PLACE_LOCATION = "NONE";
      defparam ii2057.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2058 ( .DX(nn2058), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1252_), .F3(dummy_abc_1253_) );
      defparam ii2058.CONFIG_DATA = 16'h9999;
      defparam ii2058.PLACE_LOCATION = "NONE";
      defparam ii2058.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2059 ( .DX(nn2059), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_697_) );
      defparam ii2059.CONFIG_DATA = 16'hA569;
      defparam ii2059.PLACE_LOCATION = "NONE";
      defparam ii2059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2060 ( .DX(nn2060), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_697_), .F2(nn2013), .F3(\coefcal1_divide_inst2_u110_XORCI_1|SUM_net ) );
      defparam ii2060.CONFIG_DATA = 16'hA695;
      defparam ii2060.PLACE_LOCATION = "NONE";
      defparam ii2060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2061 ( .DX(nn2061), .F0(nn2014), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_2|SUM_net ), .F3(dummy_abc_1254_) );
      defparam ii2061.CONFIG_DATA = 16'hB8B8;
      defparam ii2061.PLACE_LOCATION = "NONE";
      defparam ii2061.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2062 ( .DX(nn2062), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2061), .F2(dummy_abc_1255_), .F3(dummy_abc_1256_) );
      defparam ii2062.CONFIG_DATA = 16'h9999;
      defparam ii2062.PLACE_LOCATION = "NONE";
      defparam ii2062.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2063 ( .DX(nn2063), .F0(nn2015), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_3|SUM_net ), .F3(dummy_abc_1257_) );
      defparam ii2063.CONFIG_DATA = 16'hB8B8;
      defparam ii2063.PLACE_LOCATION = "NONE";
      defparam ii2063.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2064 ( .DX(nn2064), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2063), .F2(dummy_abc_1258_), .F3(dummy_abc_1259_) );
      defparam ii2064.CONFIG_DATA = 16'h9999;
      defparam ii2064.PLACE_LOCATION = "NONE";
      defparam ii2064.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2065 ( .DX(nn2065), .F0(nn2016), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_4|SUM_net ), .F3(dummy_abc_1260_) );
      defparam ii2065.CONFIG_DATA = 16'hB8B8;
      defparam ii2065.PLACE_LOCATION = "NONE";
      defparam ii2065.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2066 ( .DX(nn2066), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2065), .F2(dummy_abc_1261_), .F3(dummy_abc_1262_) );
      defparam ii2066.CONFIG_DATA = 16'h9999;
      defparam ii2066.PLACE_LOCATION = "NONE";
      defparam ii2066.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2067 ( .DX(nn2067), .F0(nn2017), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_5|SUM_net ), .F3(dummy_abc_1263_) );
      defparam ii2067.CONFIG_DATA = 16'hB8B8;
      defparam ii2067.PLACE_LOCATION = "NONE";
      defparam ii2067.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2068 ( .DX(nn2068), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2067), .F2(dummy_abc_1264_), .F3(dummy_abc_1265_) );
      defparam ii2068.CONFIG_DATA = 16'h9999;
      defparam ii2068.PLACE_LOCATION = "NONE";
      defparam ii2068.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2069 ( .DX(nn2069), .F0(nn2018), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_6|SUM_net ), .F3(dummy_abc_1266_) );
      defparam ii2069.CONFIG_DATA = 16'hB8B8;
      defparam ii2069.PLACE_LOCATION = "NONE";
      defparam ii2069.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2070 ( .DX(nn2070), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2069), .F2(dummy_abc_1267_), .F3(dummy_abc_1268_) );
      defparam ii2070.CONFIG_DATA = 16'h9999;
      defparam ii2070.PLACE_LOCATION = "NONE";
      defparam ii2070.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2071 ( .DX(nn2071), .F0(nn2019), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_7|SUM_net ), .F3(dummy_abc_1269_) );
      defparam ii2071.CONFIG_DATA = 16'hB8B8;
      defparam ii2071.PLACE_LOCATION = "NONE";
      defparam ii2071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2072 ( .DX(nn2072), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2071), .F2(dummy_abc_1270_), .F3(dummy_abc_1271_) );
      defparam ii2072.CONFIG_DATA = 16'h9999;
      defparam ii2072.PLACE_LOCATION = "NONE";
      defparam ii2072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2073 ( .DX(nn2073), .F0(nn2020), .F1(dummy_697_), .F2(\coefcal1_divide_inst2_u110_XORCI_8|SUM_net ), .F3(dummy_abc_1272_) );
      defparam ii2073.CONFIG_DATA = 16'hB8B8;
      defparam ii2073.PLACE_LOCATION = "NONE";
      defparam ii2073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2074 ( .DX(nn2074), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2073), .F2(dummy_abc_1273_), .F3(dummy_abc_1274_) );
      defparam ii2074.CONFIG_DATA = 16'h9999;
      defparam ii2074.PLACE_LOCATION = "NONE";
      defparam ii2074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2075 ( .DX(nn2075), .F0(dummy_678_), .F1(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ), .F2(dummy_abc_1275_), .F3(dummy_abc_1276_) );
      defparam ii2075.CONFIG_DATA = 16'h1111;
      defparam ii2075.PLACE_LOCATION = "NONE";
      defparam ii2075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2076 ( .DX(nn2076), .F0(nn1892), .F1(nn2075), .F2(dummy_697_), .F3(\coefcal1_divide_inst2_u110_XORCI_9|SUM_net ) );
      defparam ii2076.CONFIG_DATA = 16'h2A20;
      defparam ii2076.PLACE_LOCATION = "NONE";
      defparam ii2076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2077 ( .DX(nn2077), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2076), .F2(dummy_abc_1277_), .F3(dummy_abc_1278_) );
      defparam ii2077.CONFIG_DATA = 16'h9999;
      defparam ii2077.PLACE_LOCATION = "NONE";
      defparam ii2077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2078 ( .DX(nn2078), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1279_), .F2(dummy_abc_1280_), .F3(dummy_abc_1281_) );
      defparam ii2078.CONFIG_DATA = 16'h5555;
      defparam ii2078.PLACE_LOCATION = "NONE";
      defparam ii2078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2079 ( .DX(nn2079), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1282_), .F2(dummy_abc_1283_), .F3(dummy_abc_1284_) );
      defparam ii2079.CONFIG_DATA = 16'h5555;
      defparam ii2079.PLACE_LOCATION = "NONE";
      defparam ii2079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2080 ( .DX(nn2080), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1285_), .F2(dummy_abc_1286_), .F3(dummy_abc_1287_) );
      defparam ii2080.CONFIG_DATA = 16'h5555;
      defparam ii2080.PLACE_LOCATION = "NONE";
      defparam ii2080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2081 ( .DX(nn2081), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1288_), .F2(dummy_abc_1289_), .F3(dummy_abc_1290_) );
      defparam ii2081.CONFIG_DATA = 16'h5555;
      defparam ii2081.PLACE_LOCATION = "NONE";
      defparam ii2081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2082 ( .DX(nn2082), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1291_), .F2(dummy_abc_1292_), .F3(dummy_abc_1293_) );
      defparam ii2082.CONFIG_DATA = 16'h5555;
      defparam ii2082.PLACE_LOCATION = "NONE";
      defparam ii2082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2083 ( .DX(nn2083), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1294_), .F2(dummy_abc_1295_), .F3(dummy_abc_1296_) );
      defparam ii2083.CONFIG_DATA = 16'h5555;
      defparam ii2083.PLACE_LOCATION = "NONE";
      defparam ii2083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2084 ( .DX(nn2084), .F0(dummy_abc_1297_), .F1(dummy_abc_1298_), .F2(dummy_abc_1299_), .F3(dummy_abc_1300_) );
      defparam ii2084.CONFIG_DATA = 16'hFFFF;
      defparam ii2084.PLACE_LOCATION = "NONE";
      defparam ii2084.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_65_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_716_ ), 
        .DX( {nn2084, nn2083, nn2082, nn2081, nn2080, nn2079, nn2078, nn2077, 
              nn2074, nn2072, nn2070, nn2068, nn2066, nn2064, nn2062, nn2060, 
              nn2059, nn2058} ), 
        .SUM( {\coefcal1_divide_inst2_u138_XORCI_17|SUM_net , dummy_717_, 
              dummy_718_, dummy_719_, dummy_720_, dummy_721_, dummy_722_, dummy_723_, 
              dummy_724_, dummy_725_, dummy_726_, dummy_727_, dummy_728_, dummy_729_, 
              dummy_730_, dummy_731_, dummy_732_, dummy_733_} )
      );
    CS_LUT4_PRIM ii2105 ( .DX(nn2105), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_697_), .F3(dummy_abc_1301_) );
      defparam ii2105.CONFIG_DATA = 16'hA6A6;
      defparam ii2105.PLACE_LOCATION = "NONE";
      defparam ii2105.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2106 ( .DX(nn2106), .F0(dummy_697_), .F1(nn2013), .F2(\coefcal1_divide_inst2_u110_XORCI_1|SUM_net ), .F3(dummy_abc_1302_) );
      defparam ii2106.CONFIG_DATA = 16'hD8D8;
      defparam ii2106.PLACE_LOCATION = "NONE";
      defparam ii2106.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2107 ( .DX(nn2107), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1303_), .F3(dummy_abc_1304_) );
      defparam ii2107.CONFIG_DATA = 16'h9999;
      defparam ii2107.PLACE_LOCATION = "NONE";
      defparam ii2107.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2108 ( .DX(nn2108), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_697_) );
      defparam ii2108.CONFIG_DATA = 16'hA569;
      defparam ii2108.PLACE_LOCATION = "NONE";
      defparam ii2108.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2109 ( .DX(nn2109), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_697_), .F2(nn2013), .F3(\coefcal1_divide_inst2_u110_XORCI_1|SUM_net ) );
      defparam ii2109.CONFIG_DATA = 16'hA695;
      defparam ii2109.PLACE_LOCATION = "NONE";
      defparam ii2109.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2110 ( .DX(nn2110), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2061), .F2(dummy_abc_1305_), .F3(dummy_abc_1306_) );
      defparam ii2110.CONFIG_DATA = 16'h9999;
      defparam ii2110.PLACE_LOCATION = "NONE";
      defparam ii2110.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2111 ( .DX(nn2111), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2063), .F2(dummy_abc_1307_), .F3(dummy_abc_1308_) );
      defparam ii2111.CONFIG_DATA = 16'h9999;
      defparam ii2111.PLACE_LOCATION = "NONE";
      defparam ii2111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2112 ( .DX(nn2112), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2065), .F2(dummy_abc_1309_), .F3(dummy_abc_1310_) );
      defparam ii2112.CONFIG_DATA = 16'h9999;
      defparam ii2112.PLACE_LOCATION = "NONE";
      defparam ii2112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2113 ( .DX(nn2113), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2067), .F2(dummy_abc_1311_), .F3(dummy_abc_1312_) );
      defparam ii2113.CONFIG_DATA = 16'h9999;
      defparam ii2113.PLACE_LOCATION = "NONE";
      defparam ii2113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2114 ( .DX(nn2114), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2069), .F2(dummy_abc_1313_), .F3(dummy_abc_1314_) );
      defparam ii2114.CONFIG_DATA = 16'h9999;
      defparam ii2114.PLACE_LOCATION = "NONE";
      defparam ii2114.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2115 ( .DX(nn2115), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2071), .F2(dummy_abc_1315_), .F3(dummy_abc_1316_) );
      defparam ii2115.CONFIG_DATA = 16'h9999;
      defparam ii2115.PLACE_LOCATION = "NONE";
      defparam ii2115.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2116 ( .DX(nn2116), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2073), .F2(dummy_abc_1317_), .F3(dummy_abc_1318_) );
      defparam ii2116.CONFIG_DATA = 16'h9999;
      defparam ii2116.PLACE_LOCATION = "NONE";
      defparam ii2116.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2117 ( .DX(nn2117), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2076), .F2(dummy_abc_1319_), .F3(dummy_abc_1320_) );
      defparam ii2117.CONFIG_DATA = 16'h9999;
      defparam ii2117.PLACE_LOCATION = "NONE";
      defparam ii2117.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2118 ( .DX(nn2118), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1321_), .F2(dummy_abc_1322_), .F3(dummy_abc_1323_) );
      defparam ii2118.CONFIG_DATA = 16'h5555;
      defparam ii2118.PLACE_LOCATION = "NONE";
      defparam ii2118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2119 ( .DX(nn2119), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1324_), .F2(dummy_abc_1325_), .F3(dummy_abc_1326_) );
      defparam ii2119.CONFIG_DATA = 16'h5555;
      defparam ii2119.PLACE_LOCATION = "NONE";
      defparam ii2119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2120 ( .DX(nn2120), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1327_), .F2(dummy_abc_1328_), .F3(dummy_abc_1329_) );
      defparam ii2120.CONFIG_DATA = 16'h5555;
      defparam ii2120.PLACE_LOCATION = "NONE";
      defparam ii2120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2121 ( .DX(nn2121), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1330_), .F2(dummy_abc_1331_), .F3(dummy_abc_1332_) );
      defparam ii2121.CONFIG_DATA = 16'h5555;
      defparam ii2121.PLACE_LOCATION = "NONE";
      defparam ii2121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2122 ( .DX(nn2122), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1333_), .F2(dummy_abc_1334_), .F3(dummy_abc_1335_) );
      defparam ii2122.CONFIG_DATA = 16'h5555;
      defparam ii2122.PLACE_LOCATION = "NONE";
      defparam ii2122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2123 ( .DX(nn2123), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1336_), .F2(dummy_abc_1337_), .F3(dummy_abc_1338_) );
      defparam ii2123.CONFIG_DATA = 16'h5555;
      defparam ii2123.PLACE_LOCATION = "NONE";
      defparam ii2123.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_49_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn2076, nn2073, nn2071, nn2069, nn2067, nn2065, nn2063, 
              nn2061, nn2106, nn2105, \coefcal1_yDividend__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_186_ ), 
        .DX( {nn2123, nn2122, nn2121, nn2120, nn2119, nn2118, nn2117, nn2116, 
              nn2115, nn2114, nn2113, nn2112, nn2111, nn2110, nn2109, nn2108, 
              nn2107} ), 
        .SUM( {dummy_187_, \coefcal1_divide_inst2_u111_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_14|SUM_net , \coefcal1_divide_inst2_u111_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_12|SUM_net , \coefcal1_divide_inst2_u111_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_10|SUM_net , \coefcal1_divide_inst2_u111_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_8|SUM_net , \coefcal1_divide_inst2_u111_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_6|SUM_net , \coefcal1_divide_inst2_u111_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_4|SUM_net , \coefcal1_divide_inst2_u111_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_2|SUM_net , \coefcal1_divide_inst2_u111_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2143 ( .DX(nn2143), .F0(nn1892), .F1(nn2057), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_10|SUM_net ) );
      defparam ii2143.CONFIG_DATA = 16'h8A80;
      defparam ii2143.PLACE_LOCATION = "NONE";
      defparam ii2143.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2144 ( .DX(nn2144), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1339_), .F3(dummy_abc_1340_) );
      defparam ii2144.CONFIG_DATA = 16'h9999;
      defparam ii2144.PLACE_LOCATION = "NONE";
      defparam ii2144.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2145 ( .DX(nn2145), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_716_) );
      defparam ii2145.CONFIG_DATA = 16'hA569;
      defparam ii2145.PLACE_LOCATION = "NONE";
      defparam ii2145.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2146 ( .DX(nn2146), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_716_), .F2(nn2105), .F3(\coefcal1_divide_inst2_u111_XORCI_1|SUM_net ) );
      defparam ii2146.CONFIG_DATA = 16'hA695;
      defparam ii2146.PLACE_LOCATION = "NONE";
      defparam ii2146.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2147 ( .DX(nn2147), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2106), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_2|SUM_net ) );
      defparam ii2147.CONFIG_DATA = 16'h9A95;
      defparam ii2147.PLACE_LOCATION = "NONE";
      defparam ii2147.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2148 ( .DX(nn2148), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2061), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_3|SUM_net ) );
      defparam ii2148.CONFIG_DATA = 16'h9A95;
      defparam ii2148.PLACE_LOCATION = "NONE";
      defparam ii2148.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2149 ( .DX(nn2149), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2063), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_4|SUM_net ) );
      defparam ii2149.CONFIG_DATA = 16'h9A95;
      defparam ii2149.PLACE_LOCATION = "NONE";
      defparam ii2149.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2150 ( .DX(nn2150), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2065), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_5|SUM_net ) );
      defparam ii2150.CONFIG_DATA = 16'h9A95;
      defparam ii2150.PLACE_LOCATION = "NONE";
      defparam ii2150.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2151 ( .DX(nn2151), .F0(nn2067), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_6|SUM_net ), .F3(dummy_abc_1341_) );
      defparam ii2151.CONFIG_DATA = 16'hB8B8;
      defparam ii2151.PLACE_LOCATION = "NONE";
      defparam ii2151.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2152 ( .DX(nn2152), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2151), .F2(dummy_abc_1342_), .F3(dummy_abc_1343_) );
      defparam ii2152.CONFIG_DATA = 16'h9999;
      defparam ii2152.PLACE_LOCATION = "NONE";
      defparam ii2152.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2153 ( .DX(nn2153), .F0(nn2069), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_7|SUM_net ), .F3(dummy_abc_1344_) );
      defparam ii2153.CONFIG_DATA = 16'hB8B8;
      defparam ii2153.PLACE_LOCATION = "NONE";
      defparam ii2153.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2154 ( .DX(nn2154), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2153), .F2(dummy_abc_1345_), .F3(dummy_abc_1346_) );
      defparam ii2154.CONFIG_DATA = 16'h9999;
      defparam ii2154.PLACE_LOCATION = "NONE";
      defparam ii2154.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2155 ( .DX(nn2155), .F0(nn2071), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_8|SUM_net ), .F3(dummy_abc_1347_) );
      defparam ii2155.CONFIG_DATA = 16'hB8B8;
      defparam ii2155.PLACE_LOCATION = "NONE";
      defparam ii2155.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2156 ( .DX(nn2156), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2155), .F2(dummy_abc_1348_), .F3(dummy_abc_1349_) );
      defparam ii2156.CONFIG_DATA = 16'h9999;
      defparam ii2156.PLACE_LOCATION = "NONE";
      defparam ii2156.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2157 ( .DX(nn2157), .F0(nn2073), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_9|SUM_net ), .F3(dummy_abc_1350_) );
      defparam ii2157.CONFIG_DATA = 16'hB8B8;
      defparam ii2157.PLACE_LOCATION = "NONE";
      defparam ii2157.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2158 ( .DX(nn2158), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2157), .F2(dummy_abc_1351_), .F3(dummy_abc_1352_) );
      defparam ii2158.CONFIG_DATA = 16'h9999;
      defparam ii2158.PLACE_LOCATION = "NONE";
      defparam ii2158.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2159 ( .DX(nn2159), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2143), .F2(dummy_abc_1353_), .F3(dummy_abc_1354_) );
      defparam ii2159.CONFIG_DATA = 16'h9999;
      defparam ii2159.PLACE_LOCATION = "NONE";
      defparam ii2159.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2160 ( .DX(nn2160), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1355_), .F2(dummy_abc_1356_), .F3(dummy_abc_1357_) );
      defparam ii2160.CONFIG_DATA = 16'h5555;
      defparam ii2160.PLACE_LOCATION = "NONE";
      defparam ii2160.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2161 ( .DX(nn2161), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1358_), .F2(dummy_abc_1359_), .F3(dummy_abc_1360_) );
      defparam ii2161.CONFIG_DATA = 16'h5555;
      defparam ii2161.PLACE_LOCATION = "NONE";
      defparam ii2161.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2162 ( .DX(nn2162), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1361_), .F2(dummy_abc_1362_), .F3(dummy_abc_1363_) );
      defparam ii2162.CONFIG_DATA = 16'h5555;
      defparam ii2162.PLACE_LOCATION = "NONE";
      defparam ii2162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2163 ( .DX(nn2163), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1364_), .F2(dummy_abc_1365_), .F3(dummy_abc_1366_) );
      defparam ii2163.CONFIG_DATA = 16'h5555;
      defparam ii2163.PLACE_LOCATION = "NONE";
      defparam ii2163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2164 ( .DX(nn2164), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1367_), .F2(dummy_abc_1368_), .F3(dummy_abc_1369_) );
      defparam ii2164.CONFIG_DATA = 16'h5555;
      defparam ii2164.PLACE_LOCATION = "NONE";
      defparam ii2164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2165 ( .DX(nn2165), .F0(dummy_abc_1370_), .F1(dummy_abc_1371_), .F2(dummy_abc_1372_), .F3(dummy_abc_1373_) );
      defparam ii2165.CONFIG_DATA = 16'hFFFF;
      defparam ii2165.PLACE_LOCATION = "NONE";
      defparam ii2165.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_66_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_735_ ), 
        .DX( {nn2165, nn2164, nn2163, nn2162, nn2161, nn2160, nn2159, nn2158, 
              nn2156, nn2154, nn2152, nn2150, nn2149, nn2148, nn2147, nn2146, 
              nn2145, nn2144} ), 
        .SUM( {\coefcal1_divide_inst2_u140_XORCI_17|SUM_net , dummy_736_, 
              dummy_737_, dummy_738_, dummy_739_, dummy_740_, dummy_741_, dummy_742_, 
              dummy_743_, dummy_744_, dummy_745_, dummy_746_, dummy_747_, dummy_748_, 
              dummy_749_, dummy_750_, dummy_751_, dummy_752_} )
      );
    CS_LUT4_PRIM ii2186 ( .DX(nn2186), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1374_), .F3(dummy_abc_1375_) );
      defparam ii2186.CONFIG_DATA = 16'h9999;
      defparam ii2186.PLACE_LOCATION = "NONE";
      defparam ii2186.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2187 ( .DX(nn2187), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_735_) );
      defparam ii2187.CONFIG_DATA = 16'hA569;
      defparam ii2187.PLACE_LOCATION = "NONE";
      defparam ii2187.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2188 ( .DX(nn2188), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_716_), .F3(dummy_abc_1376_) );
      defparam ii2188.CONFIG_DATA = 16'hA6A6;
      defparam ii2188.PLACE_LOCATION = "NONE";
      defparam ii2188.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2189 ( .DX(nn2189), .F0(dummy_716_), .F1(nn2105), .F2(\coefcal1_divide_inst2_u111_XORCI_1|SUM_net ), .F3(dummy_abc_1377_) );
      defparam ii2189.CONFIG_DATA = 16'hD8D8;
      defparam ii2189.PLACE_LOCATION = "NONE";
      defparam ii2189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2190 ( .DX(nn2190), .F0(nn2106), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_2|SUM_net ), .F3(dummy_abc_1378_) );
      defparam ii2190.CONFIG_DATA = 16'hB8B8;
      defparam ii2190.PLACE_LOCATION = "NONE";
      defparam ii2190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2191 ( .DX(nn2191), .F0(nn2061), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_3|SUM_net ), .F3(dummy_abc_1379_) );
      defparam ii2191.CONFIG_DATA = 16'hB8B8;
      defparam ii2191.PLACE_LOCATION = "NONE";
      defparam ii2191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2192 ( .DX(nn2192), .F0(nn2063), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_4|SUM_net ), .F3(dummy_abc_1380_) );
      defparam ii2192.CONFIG_DATA = 16'hB8B8;
      defparam ii2192.PLACE_LOCATION = "NONE";
      defparam ii2192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2193 ( .DX(nn2193), .F0(nn2065), .F1(dummy_716_), .F2(\coefcal1_divide_inst2_u111_XORCI_5|SUM_net ), .F3(dummy_abc_1381_) );
      defparam ii2193.CONFIG_DATA = 16'hB8B8;
      defparam ii2193.PLACE_LOCATION = "NONE";
      defparam ii2193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2194 ( .DX(nn2194), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1382_), .F3(dummy_abc_1383_) );
      defparam ii2194.CONFIG_DATA = 16'h9999;
      defparam ii2194.PLACE_LOCATION = "NONE";
      defparam ii2194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2195 ( .DX(nn2195), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_716_) );
      defparam ii2195.CONFIG_DATA = 16'hA569;
      defparam ii2195.PLACE_LOCATION = "NONE";
      defparam ii2195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2196 ( .DX(nn2196), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_716_), .F2(nn2105), .F3(\coefcal1_divide_inst2_u111_XORCI_1|SUM_net ) );
      defparam ii2196.CONFIG_DATA = 16'hA695;
      defparam ii2196.PLACE_LOCATION = "NONE";
      defparam ii2196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2197 ( .DX(nn2197), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2106), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_2|SUM_net ) );
      defparam ii2197.CONFIG_DATA = 16'h9A95;
      defparam ii2197.PLACE_LOCATION = "NONE";
      defparam ii2197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2198 ( .DX(nn2198), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2061), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_3|SUM_net ) );
      defparam ii2198.CONFIG_DATA = 16'h9A95;
      defparam ii2198.PLACE_LOCATION = "NONE";
      defparam ii2198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2199 ( .DX(nn2199), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2063), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_4|SUM_net ) );
      defparam ii2199.CONFIG_DATA = 16'h9A95;
      defparam ii2199.PLACE_LOCATION = "NONE";
      defparam ii2199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2200 ( .DX(nn2200), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2065), .F2(dummy_716_), .F3(\coefcal1_divide_inst2_u111_XORCI_5|SUM_net ) );
      defparam ii2200.CONFIG_DATA = 16'h9A95;
      defparam ii2200.PLACE_LOCATION = "NONE";
      defparam ii2200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2201 ( .DX(nn2201), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2151), .F2(dummy_abc_1384_), .F3(dummy_abc_1385_) );
      defparam ii2201.CONFIG_DATA = 16'h9999;
      defparam ii2201.PLACE_LOCATION = "NONE";
      defparam ii2201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2202 ( .DX(nn2202), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2153), .F2(dummy_abc_1386_), .F3(dummy_abc_1387_) );
      defparam ii2202.CONFIG_DATA = 16'h9999;
      defparam ii2202.PLACE_LOCATION = "NONE";
      defparam ii2202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2203 ( .DX(nn2203), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2155), .F2(dummy_abc_1388_), .F3(dummy_abc_1389_) );
      defparam ii2203.CONFIG_DATA = 16'h9999;
      defparam ii2203.PLACE_LOCATION = "NONE";
      defparam ii2203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2204 ( .DX(nn2204), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2157), .F2(dummy_abc_1390_), .F3(dummy_abc_1391_) );
      defparam ii2204.CONFIG_DATA = 16'h9999;
      defparam ii2204.PLACE_LOCATION = "NONE";
      defparam ii2204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2205 ( .DX(nn2205), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2143), .F2(dummy_abc_1392_), .F3(dummy_abc_1393_) );
      defparam ii2205.CONFIG_DATA = 16'h9999;
      defparam ii2205.PLACE_LOCATION = "NONE";
      defparam ii2205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2206 ( .DX(nn2206), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1394_), .F2(dummy_abc_1395_), .F3(dummy_abc_1396_) );
      defparam ii2206.CONFIG_DATA = 16'h5555;
      defparam ii2206.PLACE_LOCATION = "NONE";
      defparam ii2206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2207 ( .DX(nn2207), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1397_), .F2(dummy_abc_1398_), .F3(dummy_abc_1399_) );
      defparam ii2207.CONFIG_DATA = 16'h5555;
      defparam ii2207.PLACE_LOCATION = "NONE";
      defparam ii2207.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2208 ( .DX(nn2208), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1400_), .F2(dummy_abc_1401_), .F3(dummy_abc_1402_) );
      defparam ii2208.CONFIG_DATA = 16'h5555;
      defparam ii2208.PLACE_LOCATION = "NONE";
      defparam ii2208.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2209 ( .DX(nn2209), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1403_), .F2(dummy_abc_1404_), .F3(dummy_abc_1405_) );
      defparam ii2209.CONFIG_DATA = 16'h5555;
      defparam ii2209.PLACE_LOCATION = "NONE";
      defparam ii2209.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2210 ( .DX(nn2210), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1406_), .F2(dummy_abc_1407_), .F3(dummy_abc_1408_) );
      defparam ii2210.CONFIG_DATA = 16'h5555;
      defparam ii2210.PLACE_LOCATION = "NONE";
      defparam ii2210.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_50_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2143, 
              nn2157, nn2155, nn2153, nn2151, nn2193, nn2192, nn2191, nn2190, 
              nn2189, nn2188, \coefcal1_yDividend__reg[5]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_188_ ), 
        .DX( {nn2210, nn2209, nn2208, nn2207, nn2206, nn2205, nn2204, nn2203, 
              nn2202, nn2201, nn2200, nn2199, nn2198, nn2197, nn2196, nn2195, 
              nn2194} ), 
        .SUM( {dummy_189_, \coefcal1_divide_inst2_u112_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_14|SUM_net , \coefcal1_divide_inst2_u112_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_12|SUM_net , \coefcal1_divide_inst2_u112_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_10|SUM_net , \coefcal1_divide_inst2_u112_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_8|SUM_net , \coefcal1_divide_inst2_u112_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_6|SUM_net , \coefcal1_divide_inst2_u112_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_4|SUM_net , \coefcal1_divide_inst2_u112_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_2|SUM_net , \coefcal1_divide_inst2_u112_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2230 ( .DX(nn2230), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_735_), .F2(nn2188), .F3(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ) );
      defparam ii2230.CONFIG_DATA = 16'hA695;
      defparam ii2230.PLACE_LOCATION = "NONE";
      defparam ii2230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2231 ( .DX(nn2231), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2189), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ) );
      defparam ii2231.CONFIG_DATA = 16'h9A95;
      defparam ii2231.PLACE_LOCATION = "NONE";
      defparam ii2231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2232 ( .DX(nn2232), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2190), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ) );
      defparam ii2232.CONFIG_DATA = 16'h9A95;
      defparam ii2232.PLACE_LOCATION = "NONE";
      defparam ii2232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2233 ( .DX(nn2233), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2191), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ) );
      defparam ii2233.CONFIG_DATA = 16'h9A95;
      defparam ii2233.PLACE_LOCATION = "NONE";
      defparam ii2233.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2234 ( .DX(nn2234), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2192), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ) );
      defparam ii2234.CONFIG_DATA = 16'h9A95;
      defparam ii2234.PLACE_LOCATION = "NONE";
      defparam ii2234.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2235 ( .DX(nn2235), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2193), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ) );
      defparam ii2235.CONFIG_DATA = 16'h9A95;
      defparam ii2235.PLACE_LOCATION = "NONE";
      defparam ii2235.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2236 ( .DX(nn2236), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2151), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ) );
      defparam ii2236.CONFIG_DATA = 16'h9A95;
      defparam ii2236.PLACE_LOCATION = "NONE";
      defparam ii2236.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2237 ( .DX(nn2237), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2153), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ) );
      defparam ii2237.CONFIG_DATA = 16'h9A95;
      defparam ii2237.PLACE_LOCATION = "NONE";
      defparam ii2237.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2238 ( .DX(nn2238), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2155), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ) );
      defparam ii2238.CONFIG_DATA = 16'h9A95;
      defparam ii2238.PLACE_LOCATION = "NONE";
      defparam ii2238.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2239 ( .DX(nn2239), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2157), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ) );
      defparam ii2239.CONFIG_DATA = 16'h9A95;
      defparam ii2239.PLACE_LOCATION = "NONE";
      defparam ii2239.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2240 ( .DX(nn2240), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2143), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_11|SUM_net ) );
      defparam ii2240.CONFIG_DATA = 16'h9A95;
      defparam ii2240.PLACE_LOCATION = "NONE";
      defparam ii2240.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2241 ( .DX(nn2241), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1409_), .F2(dummy_abc_1410_), .F3(dummy_abc_1411_) );
      defparam ii2241.CONFIG_DATA = 16'h5555;
      defparam ii2241.PLACE_LOCATION = "NONE";
      defparam ii2241.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2242 ( .DX(nn2242), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1412_), .F2(dummy_abc_1413_), .F3(dummy_abc_1414_) );
      defparam ii2242.CONFIG_DATA = 16'h5555;
      defparam ii2242.PLACE_LOCATION = "NONE";
      defparam ii2242.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2243 ( .DX(nn2243), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1415_), .F2(dummy_abc_1416_), .F3(dummy_abc_1417_) );
      defparam ii2243.CONFIG_DATA = 16'h5555;
      defparam ii2243.PLACE_LOCATION = "NONE";
      defparam ii2243.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2244 ( .DX(nn2244), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1418_), .F2(dummy_abc_1419_), .F3(dummy_abc_1420_) );
      defparam ii2244.CONFIG_DATA = 16'h5555;
      defparam ii2244.PLACE_LOCATION = "NONE";
      defparam ii2244.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2245 ( .DX(nn2245), .F0(dummy_abc_1421_), .F1(dummy_abc_1422_), .F2(dummy_abc_1423_), .F3(dummy_abc_1424_) );
      defparam ii2245.CONFIG_DATA = 16'hFFFF;
      defparam ii2245.PLACE_LOCATION = "NONE";
      defparam ii2245.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_67_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_754_ ), 
        .DX( {nn2245, nn2244, nn2243, nn2242, nn2241, nn2240, nn2239, nn2238, 
              nn2237, nn2236, nn2235, nn2234, nn2233, nn2232, nn2231, nn2230, 
              nn2187, nn2186} ), 
        .SUM( {\coefcal1_divide_inst2_u142_XORCI_17|SUM_net , dummy_755_, 
              dummy_756_, dummy_757_, dummy_758_, dummy_759_, dummy_760_, dummy_761_, 
              dummy_762_, dummy_763_, dummy_764_, dummy_765_, dummy_766_, dummy_767_, 
              dummy_768_, dummy_769_, dummy_770_, dummy_771_} )
      );
    CS_LUT4_PRIM ii2266 ( .DX(nn2266), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_735_), .F3(dummy_abc_1425_) );
      defparam ii2266.CONFIG_DATA = 16'hA6A6;
      defparam ii2266.PLACE_LOCATION = "NONE";
      defparam ii2266.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2267 ( .DX(nn2267), .F0(dummy_735_), .F1(nn2188), .F2(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ), .F3(dummy_abc_1426_) );
      defparam ii2267.CONFIG_DATA = 16'hD8D8;
      defparam ii2267.PLACE_LOCATION = "NONE";
      defparam ii2267.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2268 ( .DX(nn2268), .F0(nn2189), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ), .F3(dummy_abc_1427_) );
      defparam ii2268.CONFIG_DATA = 16'hB8B8;
      defparam ii2268.PLACE_LOCATION = "NONE";
      defparam ii2268.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2269 ( .DX(nn2269), .F0(nn2190), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ), .F3(dummy_abc_1428_) );
      defparam ii2269.CONFIG_DATA = 16'hB8B8;
      defparam ii2269.PLACE_LOCATION = "NONE";
      defparam ii2269.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2270 ( .DX(nn2270), .F0(nn2191), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ), .F3(dummy_abc_1429_) );
      defparam ii2270.CONFIG_DATA = 16'hB8B8;
      defparam ii2270.PLACE_LOCATION = "NONE";
      defparam ii2270.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2271 ( .DX(nn2271), .F0(nn2192), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ), .F3(dummy_abc_1430_) );
      defparam ii2271.CONFIG_DATA = 16'hB8B8;
      defparam ii2271.PLACE_LOCATION = "NONE";
      defparam ii2271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2272 ( .DX(nn2272), .F0(nn2193), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ), .F3(dummy_abc_1431_) );
      defparam ii2272.CONFIG_DATA = 16'hB8B8;
      defparam ii2272.PLACE_LOCATION = "NONE";
      defparam ii2272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2273 ( .DX(nn2273), .F0(nn2151), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ), .F3(dummy_abc_1432_) );
      defparam ii2273.CONFIG_DATA = 16'hB8B8;
      defparam ii2273.PLACE_LOCATION = "NONE";
      defparam ii2273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2274 ( .DX(nn2274), .F0(nn2153), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ), .F3(dummy_abc_1433_) );
      defparam ii2274.CONFIG_DATA = 16'hB8B8;
      defparam ii2274.PLACE_LOCATION = "NONE";
      defparam ii2274.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2275 ( .DX(nn2275), .F0(nn2155), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ), .F3(dummy_abc_1434_) );
      defparam ii2275.CONFIG_DATA = 16'hB8B8;
      defparam ii2275.PLACE_LOCATION = "NONE";
      defparam ii2275.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2276 ( .DX(nn2276), .F0(nn2157), .F1(dummy_735_), .F2(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ), .F3(dummy_abc_1435_) );
      defparam ii2276.CONFIG_DATA = 16'hB8B8;
      defparam ii2276.PLACE_LOCATION = "NONE";
      defparam ii2276.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2277 ( .DX(nn2277), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1436_), .F3(dummy_abc_1437_) );
      defparam ii2277.CONFIG_DATA = 16'h9999;
      defparam ii2277.PLACE_LOCATION = "NONE";
      defparam ii2277.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2278 ( .DX(nn2278), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_735_) );
      defparam ii2278.CONFIG_DATA = 16'hA569;
      defparam ii2278.PLACE_LOCATION = "NONE";
      defparam ii2278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2279 ( .DX(nn2279), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_735_), .F2(nn2188), .F3(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ) );
      defparam ii2279.CONFIG_DATA = 16'hA695;
      defparam ii2279.PLACE_LOCATION = "NONE";
      defparam ii2279.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2280 ( .DX(nn2280), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2189), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ) );
      defparam ii2280.CONFIG_DATA = 16'h9A95;
      defparam ii2280.PLACE_LOCATION = "NONE";
      defparam ii2280.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2281 ( .DX(nn2281), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2190), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ) );
      defparam ii2281.CONFIG_DATA = 16'h9A95;
      defparam ii2281.PLACE_LOCATION = "NONE";
      defparam ii2281.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2282 ( .DX(nn2282), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2191), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ) );
      defparam ii2282.CONFIG_DATA = 16'h9A95;
      defparam ii2282.PLACE_LOCATION = "NONE";
      defparam ii2282.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2283 ( .DX(nn2283), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2192), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ) );
      defparam ii2283.CONFIG_DATA = 16'h9A95;
      defparam ii2283.PLACE_LOCATION = "NONE";
      defparam ii2283.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2284 ( .DX(nn2284), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2193), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ) );
      defparam ii2284.CONFIG_DATA = 16'h9A95;
      defparam ii2284.PLACE_LOCATION = "NONE";
      defparam ii2284.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2285 ( .DX(nn2285), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2151), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ) );
      defparam ii2285.CONFIG_DATA = 16'h9A95;
      defparam ii2285.PLACE_LOCATION = "NONE";
      defparam ii2285.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2286 ( .DX(nn2286), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2153), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ) );
      defparam ii2286.CONFIG_DATA = 16'h9A95;
      defparam ii2286.PLACE_LOCATION = "NONE";
      defparam ii2286.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2287 ( .DX(nn2287), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2155), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ) );
      defparam ii2287.CONFIG_DATA = 16'h9A95;
      defparam ii2287.PLACE_LOCATION = "NONE";
      defparam ii2287.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2288 ( .DX(nn2288), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2157), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ) );
      defparam ii2288.CONFIG_DATA = 16'h9A95;
      defparam ii2288.PLACE_LOCATION = "NONE";
      defparam ii2288.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2289 ( .DX(nn2289), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2143), .F2(dummy_735_), .F3(\coefcal1_divide_inst2_u112_XORCI_11|SUM_net ) );
      defparam ii2289.CONFIG_DATA = 16'h9A95;
      defparam ii2289.PLACE_LOCATION = "NONE";
      defparam ii2289.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2290 ( .DX(nn2290), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1438_), .F2(dummy_abc_1439_), .F3(dummy_abc_1440_) );
      defparam ii2290.CONFIG_DATA = 16'h5555;
      defparam ii2290.PLACE_LOCATION = "NONE";
      defparam ii2290.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2291 ( .DX(nn2291), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1441_), .F2(dummy_abc_1442_), .F3(dummy_abc_1443_) );
      defparam ii2291.CONFIG_DATA = 16'h5555;
      defparam ii2291.PLACE_LOCATION = "NONE";
      defparam ii2291.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2292 ( .DX(nn2292), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1444_), .F2(dummy_abc_1445_), .F3(dummy_abc_1446_) );
      defparam ii2292.CONFIG_DATA = 16'h5555;
      defparam ii2292.PLACE_LOCATION = "NONE";
      defparam ii2292.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2293 ( .DX(nn2293), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1447_), .F2(dummy_abc_1448_), .F3(dummy_abc_1449_) );
      defparam ii2293.CONFIG_DATA = 16'h5555;
      defparam ii2293.PLACE_LOCATION = "NONE";
      defparam ii2293.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_51_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2276, 
              nn2275, nn2274, nn2273, nn2272, nn2271, nn2270, nn2269, nn2268, 
              nn2267, nn2266, \coefcal1_yDividend__reg[4]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_190_ ), 
        .DX( {nn2293, nn2292, nn2291, nn2290, nn2289, nn2288, nn2287, nn2286, 
              nn2285, nn2284, nn2283, nn2282, nn2281, nn2280, nn2279, nn2278, 
              nn2277} ), 
        .SUM( {dummy_191_, \coefcal1_divide_inst2_u113_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_14|SUM_net , \coefcal1_divide_inst2_u113_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_12|SUM_net , \coefcal1_divide_inst2_u113_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_10|SUM_net , \coefcal1_divide_inst2_u113_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_8|SUM_net , \coefcal1_divide_inst2_u113_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_6|SUM_net , \coefcal1_divide_inst2_u113_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_4|SUM_net , \coefcal1_divide_inst2_u113_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_2|SUM_net , \coefcal1_divide_inst2_u113_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2313 ( .DX(nn2313), .F0(nn2143), .F1(dummy_735_), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2313.CONFIG_DATA = 16'h8F80;
      defparam ii2313.PLACE_LOCATION = "NONE";
      defparam ii2313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2314 ( .DX(nn2314), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1450_), .F3(dummy_abc_1451_) );
      defparam ii2314.CONFIG_DATA = 16'h9999;
      defparam ii2314.PLACE_LOCATION = "NONE";
      defparam ii2314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2315 ( .DX(nn2315), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_754_) );
      defparam ii2315.CONFIG_DATA = 16'hA569;
      defparam ii2315.PLACE_LOCATION = "NONE";
      defparam ii2315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2316 ( .DX(nn2316), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_754_), .F2(nn2266), .F3(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ) );
      defparam ii2316.CONFIG_DATA = 16'hA695;
      defparam ii2316.PLACE_LOCATION = "NONE";
      defparam ii2316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2317 ( .DX(nn2317), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2267), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ) );
      defparam ii2317.CONFIG_DATA = 16'h9A95;
      defparam ii2317.PLACE_LOCATION = "NONE";
      defparam ii2317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2318 ( .DX(nn2318), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2268), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ) );
      defparam ii2318.CONFIG_DATA = 16'h9A95;
      defparam ii2318.PLACE_LOCATION = "NONE";
      defparam ii2318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2319 ( .DX(nn2319), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2269), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ) );
      defparam ii2319.CONFIG_DATA = 16'h9A95;
      defparam ii2319.PLACE_LOCATION = "NONE";
      defparam ii2319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2320 ( .DX(nn2320), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2270), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ) );
      defparam ii2320.CONFIG_DATA = 16'h9A95;
      defparam ii2320.PLACE_LOCATION = "NONE";
      defparam ii2320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2321 ( .DX(nn2321), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2271), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ) );
      defparam ii2321.CONFIG_DATA = 16'h9A95;
      defparam ii2321.PLACE_LOCATION = "NONE";
      defparam ii2321.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2322 ( .DX(nn2322), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2272), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ) );
      defparam ii2322.CONFIG_DATA = 16'h9A95;
      defparam ii2322.PLACE_LOCATION = "NONE";
      defparam ii2322.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2323 ( .DX(nn2323), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2273), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ) );
      defparam ii2323.CONFIG_DATA = 16'h9A95;
      defparam ii2323.PLACE_LOCATION = "NONE";
      defparam ii2323.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2324 ( .DX(nn2324), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2274), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ) );
      defparam ii2324.CONFIG_DATA = 16'h9A95;
      defparam ii2324.PLACE_LOCATION = "NONE";
      defparam ii2324.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2325 ( .DX(nn2325), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2275), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ) );
      defparam ii2325.CONFIG_DATA = 16'h9A95;
      defparam ii2325.PLACE_LOCATION = "NONE";
      defparam ii2325.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2326 ( .DX(nn2326), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2276), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ) );
      defparam ii2326.CONFIG_DATA = 16'h9A95;
      defparam ii2326.PLACE_LOCATION = "NONE";
      defparam ii2326.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2327 ( .DX(nn2327), .F0(nn2143), .F1(dummy_735_), .F2(dummy_abc_1452_), .F3(dummy_abc_1453_) );
      defparam ii2327.CONFIG_DATA = 16'h8888;
      defparam ii2327.PLACE_LOCATION = "NONE";
      defparam ii2327.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2328 ( .DX(nn2328), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2327), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2328.CONFIG_DATA = 16'h9095;
      defparam ii2328.PLACE_LOCATION = "NONE";
      defparam ii2328.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2329 ( .DX(nn2329), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1454_), .F2(dummy_abc_1455_), .F3(dummy_abc_1456_) );
      defparam ii2329.CONFIG_DATA = 16'h5555;
      defparam ii2329.PLACE_LOCATION = "NONE";
      defparam ii2329.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2330 ( .DX(nn2330), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1457_), .F2(dummy_abc_1458_), .F3(dummy_abc_1459_) );
      defparam ii2330.CONFIG_DATA = 16'h5555;
      defparam ii2330.PLACE_LOCATION = "NONE";
      defparam ii2330.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2331 ( .DX(nn2331), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1460_), .F2(dummy_abc_1461_), .F3(dummy_abc_1462_) );
      defparam ii2331.CONFIG_DATA = 16'h5555;
      defparam ii2331.PLACE_LOCATION = "NONE";
      defparam ii2331.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2332 ( .DX(nn2332), .F0(dummy_abc_1463_), .F1(dummy_abc_1464_), .F2(dummy_abc_1465_), .F3(dummy_abc_1466_) );
      defparam ii2332.CONFIG_DATA = 16'hFFFF;
      defparam ii2332.PLACE_LOCATION = "NONE";
      defparam ii2332.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_68_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_773_ ), 
        .DX( {nn2332, nn2331, nn2330, nn2329, nn2328, nn2326, nn2325, nn2324, 
              nn2323, nn2322, nn2321, nn2320, nn2319, nn2318, nn2317, nn2316, 
              nn2315, nn2314} ), 
        .SUM( {\coefcal1_divide_inst2_u144_XORCI_17|SUM_net , dummy_774_, 
              dummy_775_, dummy_776_, dummy_777_, dummy_778_, dummy_779_, dummy_780_, 
              dummy_781_, dummy_782_, dummy_783_, dummy_784_, dummy_785_, dummy_786_, 
              dummy_787_, dummy_788_, dummy_789_, dummy_790_} )
      );
    CS_LUT4_PRIM ii2353 ( .DX(nn2353), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_754_), .F3(dummy_abc_1467_) );
      defparam ii2353.CONFIG_DATA = 16'hA6A6;
      defparam ii2353.PLACE_LOCATION = "NONE";
      defparam ii2353.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2354 ( .DX(nn2354), .F0(dummy_754_), .F1(nn2266), .F2(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ), .F3(dummy_abc_1468_) );
      defparam ii2354.CONFIG_DATA = 16'hD8D8;
      defparam ii2354.PLACE_LOCATION = "NONE";
      defparam ii2354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2355 ( .DX(nn2355), .F0(nn2267), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ), .F3(dummy_abc_1469_) );
      defparam ii2355.CONFIG_DATA = 16'hB8B8;
      defparam ii2355.PLACE_LOCATION = "NONE";
      defparam ii2355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2356 ( .DX(nn2356), .F0(nn2268), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ), .F3(dummy_abc_1470_) );
      defparam ii2356.CONFIG_DATA = 16'hB8B8;
      defparam ii2356.PLACE_LOCATION = "NONE";
      defparam ii2356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2357 ( .DX(nn2357), .F0(nn2269), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ), .F3(dummy_abc_1471_) );
      defparam ii2357.CONFIG_DATA = 16'hB8B8;
      defparam ii2357.PLACE_LOCATION = "NONE";
      defparam ii2357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2358 ( .DX(nn2358), .F0(nn2270), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ), .F3(dummy_abc_1472_) );
      defparam ii2358.CONFIG_DATA = 16'hB8B8;
      defparam ii2358.PLACE_LOCATION = "NONE";
      defparam ii2358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2359 ( .DX(nn2359), .F0(nn2271), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ), .F3(dummy_abc_1473_) );
      defparam ii2359.CONFIG_DATA = 16'hB8B8;
      defparam ii2359.PLACE_LOCATION = "NONE";
      defparam ii2359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2360 ( .DX(nn2360), .F0(nn2272), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ), .F3(dummy_abc_1474_) );
      defparam ii2360.CONFIG_DATA = 16'hB8B8;
      defparam ii2360.PLACE_LOCATION = "NONE";
      defparam ii2360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2361 ( .DX(nn2361), .F0(nn2273), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ), .F3(dummy_abc_1475_) );
      defparam ii2361.CONFIG_DATA = 16'hB8B8;
      defparam ii2361.PLACE_LOCATION = "NONE";
      defparam ii2361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2362 ( .DX(nn2362), .F0(nn2274), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ), .F3(dummy_abc_1476_) );
      defparam ii2362.CONFIG_DATA = 16'hB8B8;
      defparam ii2362.PLACE_LOCATION = "NONE";
      defparam ii2362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2363 ( .DX(nn2363), .F0(nn2275), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ), .F3(dummy_abc_1477_) );
      defparam ii2363.CONFIG_DATA = 16'hB8B8;
      defparam ii2363.PLACE_LOCATION = "NONE";
      defparam ii2363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2364 ( .DX(nn2364), .F0(nn2276), .F1(dummy_754_), .F2(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ), .F3(dummy_abc_1478_) );
      defparam ii2364.CONFIG_DATA = 16'hB8B8;
      defparam ii2364.PLACE_LOCATION = "NONE";
      defparam ii2364.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2365 ( .DX(nn2365), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1479_), .F3(dummy_abc_1480_) );
      defparam ii2365.CONFIG_DATA = 16'h9999;
      defparam ii2365.PLACE_LOCATION = "NONE";
      defparam ii2365.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2366 ( .DX(nn2366), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_754_) );
      defparam ii2366.CONFIG_DATA = 16'hA569;
      defparam ii2366.PLACE_LOCATION = "NONE";
      defparam ii2366.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2367 ( .DX(nn2367), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_754_), .F2(nn2266), .F3(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ) );
      defparam ii2367.CONFIG_DATA = 16'hA695;
      defparam ii2367.PLACE_LOCATION = "NONE";
      defparam ii2367.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2368 ( .DX(nn2368), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2267), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ) );
      defparam ii2368.CONFIG_DATA = 16'h9A95;
      defparam ii2368.PLACE_LOCATION = "NONE";
      defparam ii2368.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2369 ( .DX(nn2369), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2268), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ) );
      defparam ii2369.CONFIG_DATA = 16'h9A95;
      defparam ii2369.PLACE_LOCATION = "NONE";
      defparam ii2369.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2370 ( .DX(nn2370), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2269), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ) );
      defparam ii2370.CONFIG_DATA = 16'h9A95;
      defparam ii2370.PLACE_LOCATION = "NONE";
      defparam ii2370.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2371 ( .DX(nn2371), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2270), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ) );
      defparam ii2371.CONFIG_DATA = 16'h9A95;
      defparam ii2371.PLACE_LOCATION = "NONE";
      defparam ii2371.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2372 ( .DX(nn2372), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2271), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ) );
      defparam ii2372.CONFIG_DATA = 16'h9A95;
      defparam ii2372.PLACE_LOCATION = "NONE";
      defparam ii2372.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2373 ( .DX(nn2373), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2272), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ) );
      defparam ii2373.CONFIG_DATA = 16'h9A95;
      defparam ii2373.PLACE_LOCATION = "NONE";
      defparam ii2373.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2374 ( .DX(nn2374), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2273), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ) );
      defparam ii2374.CONFIG_DATA = 16'h9A95;
      defparam ii2374.PLACE_LOCATION = "NONE";
      defparam ii2374.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2375 ( .DX(nn2375), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2274), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ) );
      defparam ii2375.CONFIG_DATA = 16'h9A95;
      defparam ii2375.PLACE_LOCATION = "NONE";
      defparam ii2375.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2376 ( .DX(nn2376), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2275), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ) );
      defparam ii2376.CONFIG_DATA = 16'h9A95;
      defparam ii2376.PLACE_LOCATION = "NONE";
      defparam ii2376.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2377 ( .DX(nn2377), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2276), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ) );
      defparam ii2377.CONFIG_DATA = 16'h9A95;
      defparam ii2377.PLACE_LOCATION = "NONE";
      defparam ii2377.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2378 ( .DX(nn2378), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2327), .F2(dummy_754_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2378.CONFIG_DATA = 16'h9095;
      defparam ii2378.PLACE_LOCATION = "NONE";
      defparam ii2378.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2379 ( .DX(nn2379), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1481_), .F2(dummy_abc_1482_), .F3(dummy_abc_1483_) );
      defparam ii2379.CONFIG_DATA = 16'h5555;
      defparam ii2379.PLACE_LOCATION = "NONE";
      defparam ii2379.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2380 ( .DX(nn2380), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1484_), .F2(dummy_abc_1485_), .F3(dummy_abc_1486_) );
      defparam ii2380.CONFIG_DATA = 16'h5555;
      defparam ii2380.PLACE_LOCATION = "NONE";
      defparam ii2380.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2381 ( .DX(nn2381), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1487_), .F2(dummy_abc_1488_), .F3(dummy_abc_1489_) );
      defparam ii2381.CONFIG_DATA = 16'h5555;
      defparam ii2381.PLACE_LOCATION = "NONE";
      defparam ii2381.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_52_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn2313, nn2364, nn2363, nn2362, nn2361, nn2360, nn2359, 
              nn2358, nn2357, nn2356, nn2355, nn2354, nn2353, 
              \coefcal1_yDividend__reg[3]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_192_ ), 
        .DX( {nn2381, nn2380, nn2379, nn2378, nn2377, nn2376, nn2375, nn2374, 
              nn2373, nn2372, nn2371, nn2370, nn2369, nn2368, nn2367, nn2366, 
              nn2365} ), 
        .SUM( {dummy_193_, \coefcal1_divide_inst2_u114_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_14|SUM_net , \coefcal1_divide_inst2_u114_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_12|SUM_net , \coefcal1_divide_inst2_u114_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_10|SUM_net , \coefcal1_divide_inst2_u114_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_8|SUM_net , \coefcal1_divide_inst2_u114_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_6|SUM_net , \coefcal1_divide_inst2_u114_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_4|SUM_net , \coefcal1_divide_inst2_u114_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_2|SUM_net , \coefcal1_divide_inst2_u114_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2401 ( .DX(nn2401), .F0(nn2313), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ), .F3(dummy_abc_1490_) );
      defparam ii2401.CONFIG_DATA = 16'hA8A8;
      defparam ii2401.PLACE_LOCATION = "NONE";
      defparam ii2401.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2402 ( .DX(nn2402), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1491_), .F3(dummy_abc_1492_) );
      defparam ii2402.CONFIG_DATA = 16'h9999;
      defparam ii2402.PLACE_LOCATION = "NONE";
      defparam ii2402.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2403 ( .DX(nn2403), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_773_) );
      defparam ii2403.CONFIG_DATA = 16'hA569;
      defparam ii2403.PLACE_LOCATION = "NONE";
      defparam ii2403.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2404 ( .DX(nn2404), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_773_), .F2(nn2353), .F3(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ) );
      defparam ii2404.CONFIG_DATA = 16'hA695;
      defparam ii2404.PLACE_LOCATION = "NONE";
      defparam ii2404.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2405 ( .DX(nn2405), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2354), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ) );
      defparam ii2405.CONFIG_DATA = 16'h9A95;
      defparam ii2405.PLACE_LOCATION = "NONE";
      defparam ii2405.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2406 ( .DX(nn2406), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2355), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ) );
      defparam ii2406.CONFIG_DATA = 16'h9A95;
      defparam ii2406.PLACE_LOCATION = "NONE";
      defparam ii2406.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2407 ( .DX(nn2407), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2356), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ) );
      defparam ii2407.CONFIG_DATA = 16'h9A95;
      defparam ii2407.PLACE_LOCATION = "NONE";
      defparam ii2407.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2408 ( .DX(nn2408), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2357), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ) );
      defparam ii2408.CONFIG_DATA = 16'h9A95;
      defparam ii2408.PLACE_LOCATION = "NONE";
      defparam ii2408.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2409 ( .DX(nn2409), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2358), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ) );
      defparam ii2409.CONFIG_DATA = 16'h9A95;
      defparam ii2409.PLACE_LOCATION = "NONE";
      defparam ii2409.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2410 ( .DX(nn2410), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2359), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ) );
      defparam ii2410.CONFIG_DATA = 16'h9A95;
      defparam ii2410.PLACE_LOCATION = "NONE";
      defparam ii2410.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2411 ( .DX(nn2411), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2360), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ) );
      defparam ii2411.CONFIG_DATA = 16'h9A95;
      defparam ii2411.PLACE_LOCATION = "NONE";
      defparam ii2411.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2412 ( .DX(nn2412), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2361), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ) );
      defparam ii2412.CONFIG_DATA = 16'h9A95;
      defparam ii2412.PLACE_LOCATION = "NONE";
      defparam ii2412.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2413 ( .DX(nn2413), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2362), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ) );
      defparam ii2413.CONFIG_DATA = 16'h9A95;
      defparam ii2413.PLACE_LOCATION = "NONE";
      defparam ii2413.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2414 ( .DX(nn2414), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2363), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ) );
      defparam ii2414.CONFIG_DATA = 16'h9A95;
      defparam ii2414.PLACE_LOCATION = "NONE";
      defparam ii2414.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2415 ( .DX(nn2415), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2364), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ) );
      defparam ii2415.CONFIG_DATA = 16'h9A95;
      defparam ii2415.PLACE_LOCATION = "NONE";
      defparam ii2415.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2416 ( .DX(nn2416), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2313), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ) );
      defparam ii2416.CONFIG_DATA = 16'h9995;
      defparam ii2416.PLACE_LOCATION = "NONE";
      defparam ii2416.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2417 ( .DX(nn2417), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1493_), .F2(dummy_abc_1494_), .F3(dummy_abc_1495_) );
      defparam ii2417.CONFIG_DATA = 16'h5555;
      defparam ii2417.PLACE_LOCATION = "NONE";
      defparam ii2417.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2418 ( .DX(nn2418), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1496_), .F2(dummy_abc_1497_), .F3(dummy_abc_1498_) );
      defparam ii2418.CONFIG_DATA = 16'h5555;
      defparam ii2418.PLACE_LOCATION = "NONE";
      defparam ii2418.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2419 ( .DX(nn2419), .F0(dummy_abc_1499_), .F1(dummy_abc_1500_), .F2(dummy_abc_1501_), .F3(dummy_abc_1502_) );
      defparam ii2419.CONFIG_DATA = 16'hFFFF;
      defparam ii2419.PLACE_LOCATION = "NONE";
      defparam ii2419.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_69_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_792_ ), 
        .DX( {nn2419, nn2418, nn2417, nn2416, nn2415, nn2414, nn2413, nn2412, 
              nn2411, nn2410, nn2409, nn2408, nn2407, nn2406, nn2405, nn2404, 
              nn2403, nn2402} ), 
        .SUM( {\coefcal1_divide_inst2_u146_XORCI_17|SUM_net , dummy_793_, 
              dummy_794_, dummy_795_, dummy_796_, dummy_797_, dummy_798_, dummy_799_, 
              dummy_800_, dummy_801_, dummy_802_, dummy_803_, dummy_804_, dummy_805_, 
              dummy_806_, dummy_807_, dummy_808_, dummy_809_} )
      );
    CS_LUT4_PRIM ii2440 ( .DX(nn2440), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_773_), .F3(dummy_abc_1503_) );
      defparam ii2440.CONFIG_DATA = 16'hA6A6;
      defparam ii2440.PLACE_LOCATION = "NONE";
      defparam ii2440.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2441 ( .DX(nn2441), .F0(dummy_773_), .F1(nn2353), .F2(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ), .F3(dummy_abc_1504_) );
      defparam ii2441.CONFIG_DATA = 16'hD8D8;
      defparam ii2441.PLACE_LOCATION = "NONE";
      defparam ii2441.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2442 ( .DX(nn2442), .F0(nn2354), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ), .F3(dummy_abc_1505_) );
      defparam ii2442.CONFIG_DATA = 16'hB8B8;
      defparam ii2442.PLACE_LOCATION = "NONE";
      defparam ii2442.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2443 ( .DX(nn2443), .F0(nn2355), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ), .F3(dummy_abc_1506_) );
      defparam ii2443.CONFIG_DATA = 16'hB8B8;
      defparam ii2443.PLACE_LOCATION = "NONE";
      defparam ii2443.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2444 ( .DX(nn2444), .F0(nn2356), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ), .F3(dummy_abc_1507_) );
      defparam ii2444.CONFIG_DATA = 16'hB8B8;
      defparam ii2444.PLACE_LOCATION = "NONE";
      defparam ii2444.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2445 ( .DX(nn2445), .F0(nn2357), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ), .F3(dummy_abc_1508_) );
      defparam ii2445.CONFIG_DATA = 16'hB8B8;
      defparam ii2445.PLACE_LOCATION = "NONE";
      defparam ii2445.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2446 ( .DX(nn2446), .F0(nn2358), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ), .F3(dummy_abc_1509_) );
      defparam ii2446.CONFIG_DATA = 16'hB8B8;
      defparam ii2446.PLACE_LOCATION = "NONE";
      defparam ii2446.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2447 ( .DX(nn2447), .F0(nn2359), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ), .F3(dummy_abc_1510_) );
      defparam ii2447.CONFIG_DATA = 16'hB8B8;
      defparam ii2447.PLACE_LOCATION = "NONE";
      defparam ii2447.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2448 ( .DX(nn2448), .F0(nn2360), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ), .F3(dummy_abc_1511_) );
      defparam ii2448.CONFIG_DATA = 16'hB8B8;
      defparam ii2448.PLACE_LOCATION = "NONE";
      defparam ii2448.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2449 ( .DX(nn2449), .F0(nn2361), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ), .F3(dummy_abc_1512_) );
      defparam ii2449.CONFIG_DATA = 16'hB8B8;
      defparam ii2449.PLACE_LOCATION = "NONE";
      defparam ii2449.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2450 ( .DX(nn2450), .F0(nn2362), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ), .F3(dummy_abc_1513_) );
      defparam ii2450.CONFIG_DATA = 16'hB8B8;
      defparam ii2450.PLACE_LOCATION = "NONE";
      defparam ii2450.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2451 ( .DX(nn2451), .F0(nn2363), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ), .F3(dummy_abc_1514_) );
      defparam ii2451.CONFIG_DATA = 16'hB8B8;
      defparam ii2451.PLACE_LOCATION = "NONE";
      defparam ii2451.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2452 ( .DX(nn2452), .F0(nn2364), .F1(dummy_773_), .F2(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ), .F3(dummy_abc_1515_) );
      defparam ii2452.CONFIG_DATA = 16'hB8B8;
      defparam ii2452.PLACE_LOCATION = "NONE";
      defparam ii2452.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2453 ( .DX(nn2453), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1516_), .F3(dummy_abc_1517_) );
      defparam ii2453.CONFIG_DATA = 16'h9999;
      defparam ii2453.PLACE_LOCATION = "NONE";
      defparam ii2453.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2454 ( .DX(nn2454), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_773_) );
      defparam ii2454.CONFIG_DATA = 16'hA569;
      defparam ii2454.PLACE_LOCATION = "NONE";
      defparam ii2454.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2455 ( .DX(nn2455), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_773_), .F2(nn2353), .F3(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ) );
      defparam ii2455.CONFIG_DATA = 16'hA695;
      defparam ii2455.PLACE_LOCATION = "NONE";
      defparam ii2455.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2456 ( .DX(nn2456), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2354), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ) );
      defparam ii2456.CONFIG_DATA = 16'h9A95;
      defparam ii2456.PLACE_LOCATION = "NONE";
      defparam ii2456.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2457 ( .DX(nn2457), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2355), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ) );
      defparam ii2457.CONFIG_DATA = 16'h9A95;
      defparam ii2457.PLACE_LOCATION = "NONE";
      defparam ii2457.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2458 ( .DX(nn2458), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2356), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ) );
      defparam ii2458.CONFIG_DATA = 16'h9A95;
      defparam ii2458.PLACE_LOCATION = "NONE";
      defparam ii2458.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2459 ( .DX(nn2459), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2357), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ) );
      defparam ii2459.CONFIG_DATA = 16'h9A95;
      defparam ii2459.PLACE_LOCATION = "NONE";
      defparam ii2459.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2460 ( .DX(nn2460), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2358), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ) );
      defparam ii2460.CONFIG_DATA = 16'h9A95;
      defparam ii2460.PLACE_LOCATION = "NONE";
      defparam ii2460.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2461 ( .DX(nn2461), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2359), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ) );
      defparam ii2461.CONFIG_DATA = 16'h9A95;
      defparam ii2461.PLACE_LOCATION = "NONE";
      defparam ii2461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2462 ( .DX(nn2462), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2360), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ) );
      defparam ii2462.CONFIG_DATA = 16'h9A95;
      defparam ii2462.PLACE_LOCATION = "NONE";
      defparam ii2462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2463 ( .DX(nn2463), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2361), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ) );
      defparam ii2463.CONFIG_DATA = 16'h9A95;
      defparam ii2463.PLACE_LOCATION = "NONE";
      defparam ii2463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2464 ( .DX(nn2464), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2362), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ) );
      defparam ii2464.CONFIG_DATA = 16'h9A95;
      defparam ii2464.PLACE_LOCATION = "NONE";
      defparam ii2464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2465 ( .DX(nn2465), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2363), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ) );
      defparam ii2465.CONFIG_DATA = 16'h9A95;
      defparam ii2465.PLACE_LOCATION = "NONE";
      defparam ii2465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2466 ( .DX(nn2466), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2364), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ) );
      defparam ii2466.CONFIG_DATA = 16'h9A95;
      defparam ii2466.PLACE_LOCATION = "NONE";
      defparam ii2466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2467 ( .DX(nn2467), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2313), .F2(dummy_773_), .F3(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ) );
      defparam ii2467.CONFIG_DATA = 16'h9995;
      defparam ii2467.PLACE_LOCATION = "NONE";
      defparam ii2467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2468 ( .DX(nn2468), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1518_), .F2(dummy_abc_1519_), .F3(dummy_abc_1520_) );
      defparam ii2468.CONFIG_DATA = 16'h5555;
      defparam ii2468.PLACE_LOCATION = "NONE";
      defparam ii2468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2469 ( .DX(nn2469), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1521_), .F2(dummy_abc_1522_), .F3(dummy_abc_1523_) );
      defparam ii2469.CONFIG_DATA = 16'h5555;
      defparam ii2469.PLACE_LOCATION = "NONE";
      defparam ii2469.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_53_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2401, nn2452, 
              nn2451, nn2450, nn2449, nn2448, nn2447, nn2446, nn2445, nn2444, 
              nn2443, nn2442, nn2441, nn2440, \coefcal1_yDividend__reg[2]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_194_ ), 
        .DX( {nn2469, nn2468, nn2467, nn2466, nn2465, nn2464, nn2463, nn2462, 
              nn2461, nn2460, nn2459, nn2458, nn2457, nn2456, nn2455, nn2454, 
              nn2453} ), 
        .SUM( {dummy_195_, \coefcal1_divide_inst2_u115_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_14|SUM_net , \coefcal1_divide_inst2_u115_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_12|SUM_net , \coefcal1_divide_inst2_u115_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_10|SUM_net , \coefcal1_divide_inst2_u115_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_8|SUM_net , \coefcal1_divide_inst2_u115_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_6|SUM_net , \coefcal1_divide_inst2_u115_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_4|SUM_net , \coefcal1_divide_inst2_u115_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_2|SUM_net , \coefcal1_divide_inst2_u115_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2489 ( .DX(nn2489), .F0(nn2401), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_14|SUM_net ), .F3(dummy_abc_1524_) );
      defparam ii2489.CONFIG_DATA = 16'hB8B8;
      defparam ii2489.PLACE_LOCATION = "NONE";
      defparam ii2489.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2490 ( .DX(nn2490), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1525_), .F3(dummy_abc_1526_) );
      defparam ii2490.CONFIG_DATA = 16'h9999;
      defparam ii2490.PLACE_LOCATION = "NONE";
      defparam ii2490.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2491 ( .DX(nn2491), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_792_) );
      defparam ii2491.CONFIG_DATA = 16'hA569;
      defparam ii2491.PLACE_LOCATION = "NONE";
      defparam ii2491.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2492 ( .DX(nn2492), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_792_), .F2(nn2440), .F3(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ) );
      defparam ii2492.CONFIG_DATA = 16'hA695;
      defparam ii2492.PLACE_LOCATION = "NONE";
      defparam ii2492.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2493 ( .DX(nn2493), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2441), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ) );
      defparam ii2493.CONFIG_DATA = 16'h9A95;
      defparam ii2493.PLACE_LOCATION = "NONE";
      defparam ii2493.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2494 ( .DX(nn2494), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2442), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ) );
      defparam ii2494.CONFIG_DATA = 16'h9A95;
      defparam ii2494.PLACE_LOCATION = "NONE";
      defparam ii2494.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2495 ( .DX(nn2495), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2443), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ) );
      defparam ii2495.CONFIG_DATA = 16'h9A95;
      defparam ii2495.PLACE_LOCATION = "NONE";
      defparam ii2495.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2496 ( .DX(nn2496), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2444), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ) );
      defparam ii2496.CONFIG_DATA = 16'h9A95;
      defparam ii2496.PLACE_LOCATION = "NONE";
      defparam ii2496.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2497 ( .DX(nn2497), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2445), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ) );
      defparam ii2497.CONFIG_DATA = 16'h9A95;
      defparam ii2497.PLACE_LOCATION = "NONE";
      defparam ii2497.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2498 ( .DX(nn2498), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2446), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ) );
      defparam ii2498.CONFIG_DATA = 16'h9A95;
      defparam ii2498.PLACE_LOCATION = "NONE";
      defparam ii2498.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2499 ( .DX(nn2499), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2447), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ) );
      defparam ii2499.CONFIG_DATA = 16'h9A95;
      defparam ii2499.PLACE_LOCATION = "NONE";
      defparam ii2499.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2500 ( .DX(nn2500), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2448), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ) );
      defparam ii2500.CONFIG_DATA = 16'h9A95;
      defparam ii2500.PLACE_LOCATION = "NONE";
      defparam ii2500.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2501 ( .DX(nn2501), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2449), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_10|SUM_net ) );
      defparam ii2501.CONFIG_DATA = 16'h9A95;
      defparam ii2501.PLACE_LOCATION = "NONE";
      defparam ii2501.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2502 ( .DX(nn2502), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2450), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_11|SUM_net ) );
      defparam ii2502.CONFIG_DATA = 16'h9A95;
      defparam ii2502.PLACE_LOCATION = "NONE";
      defparam ii2502.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2503 ( .DX(nn2503), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2451), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_12|SUM_net ) );
      defparam ii2503.CONFIG_DATA = 16'h9A95;
      defparam ii2503.PLACE_LOCATION = "NONE";
      defparam ii2503.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2504 ( .DX(nn2504), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2452), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_13|SUM_net ) );
      defparam ii2504.CONFIG_DATA = 16'h9A95;
      defparam ii2504.PLACE_LOCATION = "NONE";
      defparam ii2504.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2505 ( .DX(nn2505), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2401), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_14|SUM_net ) );
      defparam ii2505.CONFIG_DATA = 16'h9A95;
      defparam ii2505.PLACE_LOCATION = "NONE";
      defparam ii2505.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2506 ( .DX(nn2506), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1527_), .F2(dummy_abc_1528_), .F3(dummy_abc_1529_) );
      defparam ii2506.CONFIG_DATA = 16'h5555;
      defparam ii2506.PLACE_LOCATION = "NONE";
      defparam ii2506.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2507 ( .DX(nn2507), .F0(dummy_abc_1530_), .F1(dummy_abc_1531_), .F2(dummy_abc_1532_), .F3(dummy_abc_1533_) );
      defparam ii2507.CONFIG_DATA = 16'hFFFF;
      defparam ii2507.PLACE_LOCATION = "NONE";
      defparam ii2507.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_70_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_811_ ), 
        .DX( {nn2507, nn2506, nn2505, nn2504, nn2503, nn2502, nn2501, nn2500, 
              nn2499, nn2498, nn2497, nn2496, nn2495, nn2494, nn2493, nn2492, 
              nn2491, nn2490} ), 
        .SUM( {\coefcal1_divide_inst2_u148_XORCI_17|SUM_net , dummy_812_, 
              dummy_813_, dummy_814_, dummy_815_, dummy_816_, dummy_817_, dummy_818_, 
              dummy_819_, dummy_820_, dummy_821_, dummy_822_, dummy_823_, dummy_824_, 
              dummy_825_, dummy_826_, dummy_827_, dummy_828_} )
      );
    CS_LUT4_PRIM ii2528 ( .DX(nn2528), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_792_), .F3(dummy_abc_1534_) );
      defparam ii2528.CONFIG_DATA = 16'hA6A6;
      defparam ii2528.PLACE_LOCATION = "NONE";
      defparam ii2528.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2529 ( .DX(nn2529), .F0(dummy_792_), .F1(nn2440), .F2(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ), .F3(dummy_abc_1535_) );
      defparam ii2529.CONFIG_DATA = 16'hD8D8;
      defparam ii2529.PLACE_LOCATION = "NONE";
      defparam ii2529.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2530 ( .DX(nn2530), .F0(nn2441), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ), .F3(dummy_abc_1536_) );
      defparam ii2530.CONFIG_DATA = 16'hB8B8;
      defparam ii2530.PLACE_LOCATION = "NONE";
      defparam ii2530.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2531 ( .DX(nn2531), .F0(nn2442), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ), .F3(dummy_abc_1537_) );
      defparam ii2531.CONFIG_DATA = 16'hB8B8;
      defparam ii2531.PLACE_LOCATION = "NONE";
      defparam ii2531.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2532 ( .DX(nn2532), .F0(nn2443), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ), .F3(dummy_abc_1538_) );
      defparam ii2532.CONFIG_DATA = 16'hB8B8;
      defparam ii2532.PLACE_LOCATION = "NONE";
      defparam ii2532.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2533 ( .DX(nn2533), .F0(nn2444), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ), .F3(dummy_abc_1539_) );
      defparam ii2533.CONFIG_DATA = 16'hB8B8;
      defparam ii2533.PLACE_LOCATION = "NONE";
      defparam ii2533.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2534 ( .DX(nn2534), .F0(nn2445), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ), .F3(dummy_abc_1540_) );
      defparam ii2534.CONFIG_DATA = 16'hB8B8;
      defparam ii2534.PLACE_LOCATION = "NONE";
      defparam ii2534.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2535 ( .DX(nn2535), .F0(nn2446), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ), .F3(dummy_abc_1541_) );
      defparam ii2535.CONFIG_DATA = 16'hB8B8;
      defparam ii2535.PLACE_LOCATION = "NONE";
      defparam ii2535.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2536 ( .DX(nn2536), .F0(nn2447), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ), .F3(dummy_abc_1542_) );
      defparam ii2536.CONFIG_DATA = 16'hB8B8;
      defparam ii2536.PLACE_LOCATION = "NONE";
      defparam ii2536.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2537 ( .DX(nn2537), .F0(nn2448), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ), .F3(dummy_abc_1543_) );
      defparam ii2537.CONFIG_DATA = 16'hB8B8;
      defparam ii2537.PLACE_LOCATION = "NONE";
      defparam ii2537.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2538 ( .DX(nn2538), .F0(nn2449), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_10|SUM_net ), .F3(dummy_abc_1544_) );
      defparam ii2538.CONFIG_DATA = 16'hB8B8;
      defparam ii2538.PLACE_LOCATION = "NONE";
      defparam ii2538.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2539 ( .DX(nn2539), .F0(nn2450), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_11|SUM_net ), .F3(dummy_abc_1545_) );
      defparam ii2539.CONFIG_DATA = 16'hB8B8;
      defparam ii2539.PLACE_LOCATION = "NONE";
      defparam ii2539.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2540 ( .DX(nn2540), .F0(nn2451), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_12|SUM_net ), .F3(dummy_abc_1546_) );
      defparam ii2540.CONFIG_DATA = 16'hB8B8;
      defparam ii2540.PLACE_LOCATION = "NONE";
      defparam ii2540.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2541 ( .DX(nn2541), .F0(nn2452), .F1(dummy_792_), .F2(\coefcal1_divide_inst2_u115_XORCI_13|SUM_net ), .F3(dummy_abc_1547_) );
      defparam ii2541.CONFIG_DATA = 16'hB8B8;
      defparam ii2541.PLACE_LOCATION = "NONE";
      defparam ii2541.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2542 ( .DX(nn2542), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1548_), .F3(dummy_abc_1549_) );
      defparam ii2542.CONFIG_DATA = 16'h9999;
      defparam ii2542.PLACE_LOCATION = "NONE";
      defparam ii2542.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2543 ( .DX(nn2543), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_792_) );
      defparam ii2543.CONFIG_DATA = 16'hA569;
      defparam ii2543.PLACE_LOCATION = "NONE";
      defparam ii2543.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2544 ( .DX(nn2544), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_792_), .F2(nn2440), .F3(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ) );
      defparam ii2544.CONFIG_DATA = 16'hA695;
      defparam ii2544.PLACE_LOCATION = "NONE";
      defparam ii2544.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2545 ( .DX(nn2545), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2441), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ) );
      defparam ii2545.CONFIG_DATA = 16'h9A95;
      defparam ii2545.PLACE_LOCATION = "NONE";
      defparam ii2545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2546 ( .DX(nn2546), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2442), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ) );
      defparam ii2546.CONFIG_DATA = 16'h9A95;
      defparam ii2546.PLACE_LOCATION = "NONE";
      defparam ii2546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2547 ( .DX(nn2547), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2443), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ) );
      defparam ii2547.CONFIG_DATA = 16'h9A95;
      defparam ii2547.PLACE_LOCATION = "NONE";
      defparam ii2547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2548 ( .DX(nn2548), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2444), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ) );
      defparam ii2548.CONFIG_DATA = 16'h9A95;
      defparam ii2548.PLACE_LOCATION = "NONE";
      defparam ii2548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2549 ( .DX(nn2549), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2445), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ) );
      defparam ii2549.CONFIG_DATA = 16'h9A95;
      defparam ii2549.PLACE_LOCATION = "NONE";
      defparam ii2549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2550 ( .DX(nn2550), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2446), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ) );
      defparam ii2550.CONFIG_DATA = 16'h9A95;
      defparam ii2550.PLACE_LOCATION = "NONE";
      defparam ii2550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2551 ( .DX(nn2551), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2447), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ) );
      defparam ii2551.CONFIG_DATA = 16'h9A95;
      defparam ii2551.PLACE_LOCATION = "NONE";
      defparam ii2551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2552 ( .DX(nn2552), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2448), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ) );
      defparam ii2552.CONFIG_DATA = 16'h9A95;
      defparam ii2552.PLACE_LOCATION = "NONE";
      defparam ii2552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2553 ( .DX(nn2553), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2449), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_10|SUM_net ) );
      defparam ii2553.CONFIG_DATA = 16'h9A95;
      defparam ii2553.PLACE_LOCATION = "NONE";
      defparam ii2553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2554 ( .DX(nn2554), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2450), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_11|SUM_net ) );
      defparam ii2554.CONFIG_DATA = 16'h9A95;
      defparam ii2554.PLACE_LOCATION = "NONE";
      defparam ii2554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2555 ( .DX(nn2555), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2451), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_12|SUM_net ) );
      defparam ii2555.CONFIG_DATA = 16'h9A95;
      defparam ii2555.PLACE_LOCATION = "NONE";
      defparam ii2555.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2556 ( .DX(nn2556), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2452), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_13|SUM_net ) );
      defparam ii2556.CONFIG_DATA = 16'h9A95;
      defparam ii2556.PLACE_LOCATION = "NONE";
      defparam ii2556.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2557 ( .DX(nn2557), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2401), .F2(dummy_792_), .F3(\coefcal1_divide_inst2_u115_XORCI_14|SUM_net ) );
      defparam ii2557.CONFIG_DATA = 16'h9A95;
      defparam ii2557.PLACE_LOCATION = "NONE";
      defparam ii2557.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2558 ( .DX(nn2558), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1550_), .F2(dummy_abc_1551_), .F3(dummy_abc_1552_) );
      defparam ii2558.CONFIG_DATA = 16'h5555;
      defparam ii2558.PLACE_LOCATION = "NONE";
      defparam ii2558.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_54_ ( 
        .CA( {a_acc_en_cal1_u134_mac, nn2489, nn2541, nn2540, nn2539, nn2538, 
              nn2537, nn2536, nn2535, nn2534, nn2533, nn2532, nn2531, nn2530, 
              nn2529, nn2528, \coefcal1_yDividend__reg[1]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_196_ ), 
        .DX( {nn2558, nn2557, nn2556, nn2555, nn2554, nn2553, nn2552, nn2551, 
              nn2550, nn2549, nn2548, nn2547, nn2546, nn2545, nn2544, nn2543, 
              nn2542} ), 
        .SUM( {dummy_197_, \coefcal1_divide_inst2_u116_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_14|SUM_net , \coefcal1_divide_inst2_u116_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_12|SUM_net , \coefcal1_divide_inst2_u116_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_10|SUM_net , \coefcal1_divide_inst2_u116_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_8|SUM_net , \coefcal1_divide_inst2_u116_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_6|SUM_net , \coefcal1_divide_inst2_u116_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_4|SUM_net , \coefcal1_divide_inst2_u116_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_2|SUM_net , \coefcal1_divide_inst2_u116_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2578 ( .DX(nn2578), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(nn2489), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_15|SUM_net ) );
      defparam ii2578.CONFIG_DATA = 16'h8A80;
      defparam ii2578.PLACE_LOCATION = "NONE";
      defparam ii2578.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2579 ( .DX(nn2579), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[16]|Q_net ), .F2(nn2578), .F3(dummy_abc_1553_) );
      defparam ii2579.CONFIG_DATA = 16'hF1F1;
      defparam ii2579.PLACE_LOCATION = "NONE";
      defparam ii2579.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2580 ( .DX(nn2580), .F0(dummy_abc_1554_), .F1(dummy_abc_1555_), .F2(dummy_abc_1556_), .F3(dummy_abc_1557_) );
      defparam ii2580.CONFIG_DATA = 16'hFFFF;
      defparam ii2580.PLACE_LOCATION = "NONE";
      defparam ii2580.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_55_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDividend__reg[16]|Q_net , 
              \coefcal1_yDividend__reg[15]|Q_net , \coefcal1_yDividend__reg[14]|Q_net , 
              \coefcal1_yDividend__reg[13]|Q_net , \coefcal1_yDividend__reg[12]|Q_net , 
              \coefcal1_yDividend__reg[11]|Q_net , \coefcal1_yDividend__reg[10]|Q_net , 
              \coefcal1_yDividend__reg[9]|Q_net , \coefcal1_yDividend__reg[8]|Q_net , 
              \coefcal1_yDividend__reg[7]|Q_net , \coefcal1_yDividend__reg[6]|Q_net , 
              \coefcal1_yDividend__reg[5]|Q_net , \coefcal1_yDividend__reg[4]|Q_net , 
              \coefcal1_yDividend__reg[3]|Q_net , \coefcal1_yDividend__reg[2]|Q_net , 
              \coefcal1_yDividend__reg[1]|Q_net , \coefcal1_yDividend__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_526_ ), 
        .DX( {nn2580, nn2579, nn1347, nn1346, nn1345, nn1344, nn1343, nn1342, 
              nn1341, nn1340, nn1339, nn1338, nn1337, nn1336, nn1335, nn1334, 
              nn1333, nn1332} ), 
        .SUM( {\coefcal1_divide_inst2_u118_XORCI_17|SUM_net , dummy_527_, 
              dummy_528_, dummy_529_, dummy_530_, dummy_531_, dummy_532_, dummy_533_, 
              dummy_534_, dummy_535_, dummy_536_, dummy_537_, dummy_538_, dummy_539_, 
              dummy_540_, dummy_541_, dummy_542_, dummy_543_} )
      );
    CS_LUT4_PRIM ii2601 ( .DX(nn2601), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1558_), .F3(dummy_abc_1559_) );
      defparam ii2601.CONFIG_DATA = 16'h9999;
      defparam ii2601.PLACE_LOCATION = "NONE";
      defparam ii2601.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2602 ( .DX(nn2602), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_811_) );
      defparam ii2602.CONFIG_DATA = 16'hA569;
      defparam ii2602.PLACE_LOCATION = "NONE";
      defparam ii2602.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2603 ( .DX(nn2603), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_811_), .F2(nn2528), .F3(\coefcal1_divide_inst2_u116_XORCI_1|SUM_net ) );
      defparam ii2603.CONFIG_DATA = 16'hA695;
      defparam ii2603.PLACE_LOCATION = "NONE";
      defparam ii2603.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2604 ( .DX(nn2604), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2529), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_2|SUM_net ) );
      defparam ii2604.CONFIG_DATA = 16'h9A95;
      defparam ii2604.PLACE_LOCATION = "NONE";
      defparam ii2604.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2605 ( .DX(nn2605), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2530), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_3|SUM_net ) );
      defparam ii2605.CONFIG_DATA = 16'h9A95;
      defparam ii2605.PLACE_LOCATION = "NONE";
      defparam ii2605.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2606 ( .DX(nn2606), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2531), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_4|SUM_net ) );
      defparam ii2606.CONFIG_DATA = 16'h9A95;
      defparam ii2606.PLACE_LOCATION = "NONE";
      defparam ii2606.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2607 ( .DX(nn2607), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2532), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_5|SUM_net ) );
      defparam ii2607.CONFIG_DATA = 16'h9A95;
      defparam ii2607.PLACE_LOCATION = "NONE";
      defparam ii2607.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2608 ( .DX(nn2608), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2533), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_6|SUM_net ) );
      defparam ii2608.CONFIG_DATA = 16'h9A95;
      defparam ii2608.PLACE_LOCATION = "NONE";
      defparam ii2608.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2609 ( .DX(nn2609), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2534), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_7|SUM_net ) );
      defparam ii2609.CONFIG_DATA = 16'h9A95;
      defparam ii2609.PLACE_LOCATION = "NONE";
      defparam ii2609.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2610 ( .DX(nn2610), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2535), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_8|SUM_net ) );
      defparam ii2610.CONFIG_DATA = 16'h9A95;
      defparam ii2610.PLACE_LOCATION = "NONE";
      defparam ii2610.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2611 ( .DX(nn2611), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2536), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_9|SUM_net ) );
      defparam ii2611.CONFIG_DATA = 16'h9A95;
      defparam ii2611.PLACE_LOCATION = "NONE";
      defparam ii2611.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2612 ( .DX(nn2612), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2537), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_10|SUM_net ) );
      defparam ii2612.CONFIG_DATA = 16'h9A95;
      defparam ii2612.PLACE_LOCATION = "NONE";
      defparam ii2612.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2613 ( .DX(nn2613), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2538), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_11|SUM_net ) );
      defparam ii2613.CONFIG_DATA = 16'h9A95;
      defparam ii2613.PLACE_LOCATION = "NONE";
      defparam ii2613.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2614 ( .DX(nn2614), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2539), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_12|SUM_net ) );
      defparam ii2614.CONFIG_DATA = 16'h9A95;
      defparam ii2614.PLACE_LOCATION = "NONE";
      defparam ii2614.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2615 ( .DX(nn2615), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2540), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_13|SUM_net ) );
      defparam ii2615.CONFIG_DATA = 16'h9A95;
      defparam ii2615.PLACE_LOCATION = "NONE";
      defparam ii2615.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2616 ( .DX(nn2616), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2541), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_14|SUM_net ) );
      defparam ii2616.CONFIG_DATA = 16'h9A95;
      defparam ii2616.PLACE_LOCATION = "NONE";
      defparam ii2616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2617 ( .DX(nn2617), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(nn2489), .F2(dummy_811_), .F3(\coefcal1_divide_inst2_u116_XORCI_15|SUM_net ) );
      defparam ii2617.CONFIG_DATA = 16'h9A95;
      defparam ii2617.PLACE_LOCATION = "NONE";
      defparam ii2617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2618 ( .DX(nn2618), .F0(dummy_abc_1560_), .F1(dummy_abc_1561_), .F2(dummy_abc_1562_), .F3(dummy_abc_1563_) );
      defparam ii2618.CONFIG_DATA = 16'hFFFF;
      defparam ii2618.PLACE_LOCATION = "NONE";
      defparam ii2618.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_71_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_830_ ), 
        .DX( {nn2618, nn2617, nn2616, nn2615, nn2614, nn2613, nn2612, nn2611, 
              nn2610, nn2609, nn2608, nn2607, nn2606, nn2605, nn2604, nn2603, 
              nn2602, nn2601} ), 
        .SUM( {\coefcal1_divide_inst2_u150_XORCI_17|SUM_net , dummy_831_, 
              dummy_832_, dummy_833_, dummy_834_, dummy_835_, dummy_836_, dummy_837_, 
              dummy_838_, dummy_839_, dummy_840_, dummy_841_, dummy_842_, dummy_843_, 
              dummy_844_, dummy_845_, dummy_846_, dummy_847_} )
      );
    CS_LUT4_PRIM ii2639 ( .DX(nn2639), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[7]|Q_net ), .F2(\coefcal1_yDivisor__reg[8]|Q_net ), .F3(\coefcal1_yDivisor__reg[9]|Q_net ) );
      defparam ii2639.CONFIG_DATA = 16'h0001;
      defparam ii2639.PLACE_LOCATION = "NONE";
      defparam ii2639.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2640 ( .DX(nn2640), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(\coefcal1_yDivisor__reg[5]|Q_net ), .F3(nn2639) );
      defparam ii2640.CONFIG_DATA = 16'h0100;
      defparam ii2640.PLACE_LOCATION = "NONE";
      defparam ii2640.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2641 ( .DX(nn2641), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[15]|Q_net ), .F2(\coefcal1_yDivisor__reg[16]|Q_net ), .F3(\coefcal1_yDivisor__reg[1]|Q_net ) );
      defparam ii2641.CONFIG_DATA = 16'h0001;
      defparam ii2641.PLACE_LOCATION = "NONE";
      defparam ii2641.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2642 ( .DX(nn2642), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[11]|Q_net ), .F2(\coefcal1_yDivisor__reg[12]|Q_net ), .F3(nn2641) );
      defparam ii2642.CONFIG_DATA = 16'h0100;
      defparam ii2642.PLACE_LOCATION = "NONE";
      defparam ii2642.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2643 ( .DX(nn2643), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[4]|Q_net ), .F2(nn2640), .F3(nn2642) );
      defparam ii2643.CONFIG_DATA = 16'h1000;
      defparam ii2643.PLACE_LOCATION = "NONE";
      defparam ii2643.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2644 ( .DX(nn2644), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_830_), .F3(nn2643) );
      defparam ii2644.CONFIG_DATA = 16'h77F0;
      defparam ii2644.PLACE_LOCATION = "NONE";
      defparam ii2644.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2645 ( .DX(nn2645), .F0(rst), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_526_), .F3(nn2644) );
      defparam ii2645.CONFIG_DATA = 16'h3363;
      defparam ii2645.PLACE_LOCATION = "NONE";
      defparam ii2645.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2646 ( .DX(nn2646), .F0(rst), .F1(dummy_526_), .F2(nn2644), .F3(dummy_abc_1564_) );
      defparam ii2646.CONFIG_DATA = 16'hFBFB;
      defparam ii2646.PLACE_LOCATION = "NONE";
      defparam ii2646.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2647 ( .DX(nn2647), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_811_), .F3(nn2643) );
      defparam ii2647.CONFIG_DATA = 16'h77F0;
      defparam ii2647.PLACE_LOCATION = "NONE";
      defparam ii2647.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2648 ( .DX(nn2648), .F0(rst), .F1(dummy_526_), .F2(nn2647), .F3(dummy_abc_1565_) );
      defparam ii2648.CONFIG_DATA = 16'h0404;
      defparam ii2648.PLACE_LOCATION = "NONE";
      defparam ii2648.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2649 ( .DX(nn2649), .F0(rst), .F1(\coefcal1_yDividend__reg[2]|Q_net ), .F2(\coefcal1_yDivisor__reg[0]|Q_net ), .F3(nn2643) );
      defparam ii2649.CONFIG_DATA = 16'h4055;
      defparam ii2649.PLACE_LOCATION = "NONE";
      defparam ii2649.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2650 ( .DX(nn2650), .F0(dummy_792_), .F1(dummy_526_), .F2(nn2643), .F3(nn2649) );
      defparam ii2650.CONFIG_DATA = 16'hC400;
      defparam ii2650.PLACE_LOCATION = "NONE";
      defparam ii2650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2651 ( .DX(nn2651), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_773_), .F3(nn2643) );
      defparam ii2651.CONFIG_DATA = 16'h880F;
      defparam ii2651.PLACE_LOCATION = "NONE";
      defparam ii2651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2652 ( .DX(nn2652), .F0(rst), .F1(dummy_526_), .F2(nn2651), .F3(dummy_abc_1566_) );
      defparam ii2652.CONFIG_DATA = 16'h4040;
      defparam ii2652.PLACE_LOCATION = "NONE";
      defparam ii2652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2653 ( .DX(nn2653), .F0(rst), .F1(\coefcal1_yDividend__reg[4]|Q_net ), .F2(\coefcal1_yDivisor__reg[0]|Q_net ), .F3(nn2643) );
      defparam ii2653.CONFIG_DATA = 16'h4055;
      defparam ii2653.PLACE_LOCATION = "NONE";
      defparam ii2653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2654 ( .DX(nn2654), .F0(dummy_754_), .F1(dummy_526_), .F2(nn2643), .F3(nn2653) );
      defparam ii2654.CONFIG_DATA = 16'hC400;
      defparam ii2654.PLACE_LOCATION = "NONE";
      defparam ii2654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2655 ( .DX(nn2655), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_735_), .F3(nn2643) );
      defparam ii2655.CONFIG_DATA = 16'h880F;
      defparam ii2655.PLACE_LOCATION = "NONE";
      defparam ii2655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2656 ( .DX(nn2656), .F0(rst), .F1(dummy_526_), .F2(nn2655), .F3(dummy_abc_1567_) );
      defparam ii2656.CONFIG_DATA = 16'h4040;
      defparam ii2656.PLACE_LOCATION = "NONE";
      defparam ii2656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2657 ( .DX(nn2657), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_716_), .F3(nn2643) );
      defparam ii2657.CONFIG_DATA = 16'h77F0;
      defparam ii2657.PLACE_LOCATION = "NONE";
      defparam ii2657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2658 ( .DX(nn2658), .F0(rst), .F1(dummy_526_), .F2(nn2657), .F3(dummy_abc_1568_) );
      defparam ii2658.CONFIG_DATA = 16'h0404;
      defparam ii2658.PLACE_LOCATION = "NONE";
      defparam ii2658.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2659 ( .DX(nn2659), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_697_), .F3(nn2643) );
      defparam ii2659.CONFIG_DATA = 16'h77F0;
      defparam ii2659.PLACE_LOCATION = "NONE";
      defparam ii2659.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2660 ( .DX(nn2660), .F0(rst), .F1(dummy_526_), .F2(nn2659), .F3(dummy_abc_1569_) );
      defparam ii2660.CONFIG_DATA = 16'h0404;
      defparam ii2660.PLACE_LOCATION = "NONE";
      defparam ii2660.PCK_LOCATION = "NONE";
    scaler_ipc_adder_8 carry_8_74_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_dinxy_cen_cal1_u134_mac} ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_887_ ), 
        .DX( {nn2660, nn2658, nn2656, nn2654, nn2652, nn2650, nn2648, nn2646} ), 
        .SUM( {\coefcal1_u62_XORCI_7|SUM_net , \coefcal1_u62_XORCI_6|SUM_net , 
              \coefcal1_u62_XORCI_5|SUM_net , \coefcal1_u62_XORCI_4|SUM_net , 
              \coefcal1_u62_XORCI_3|SUM_net , \coefcal1_u62_XORCI_2|SUM_net , 
              \coefcal1_u62_XORCI_1|SUM_net , \coefcal1_u62_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2671 ( .DX(nn2671), .F0(\cal1_v__reg[1]|Q_net ), .F1(\coefcal1_u62_XORCI_1|SUM_net ), .F2(dummy_abc_1570_), .F3(dummy_abc_1571_) );
      defparam ii2671.CONFIG_DATA = 16'h6666;
      defparam ii2671.PLACE_LOCATION = "NONE";
      defparam ii2671.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2672 ( .DX(nn2672), .F0(\cal1_v__reg[2]|Q_net ), .F1(\coefcal1_u62_XORCI_2|SUM_net ), .F2(dummy_abc_1572_), .F3(dummy_abc_1573_) );
      defparam ii2672.CONFIG_DATA = 16'h6666;
      defparam ii2672.PLACE_LOCATION = "NONE";
      defparam ii2672.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2673 ( .DX(nn2673), .F0(\cal1_v__reg[3]|Q_net ), .F1(\coefcal1_u62_XORCI_3|SUM_net ), .F2(dummy_abc_1574_), .F3(dummy_abc_1575_) );
      defparam ii2673.CONFIG_DATA = 16'h6666;
      defparam ii2673.PLACE_LOCATION = "NONE";
      defparam ii2673.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2674 ( .DX(nn2674), .F0(\cal1_v__reg[4]|Q_net ), .F1(\coefcal1_u62_XORCI_4|SUM_net ), .F2(dummy_abc_1576_), .F3(dummy_abc_1577_) );
      defparam ii2674.CONFIG_DATA = 16'h6666;
      defparam ii2674.PLACE_LOCATION = "NONE";
      defparam ii2674.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2675 ( .DX(nn2675), .F0(\cal1_v__reg[5]|Q_net ), .F1(\coefcal1_u62_XORCI_5|SUM_net ), .F2(dummy_abc_1578_), .F3(dummy_abc_1579_) );
      defparam ii2675.CONFIG_DATA = 16'h6666;
      defparam ii2675.PLACE_LOCATION = "NONE";
      defparam ii2675.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2676 ( .DX(nn2676), .F0(\cal1_v__reg[6]|Q_net ), .F1(\coefcal1_u62_XORCI_6|SUM_net ), .F2(dummy_abc_1580_), .F3(dummy_abc_1581_) );
      defparam ii2676.CONFIG_DATA = 16'h6666;
      defparam ii2676.PLACE_LOCATION = "NONE";
      defparam ii2676.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2677 ( .DX(nn2677), .F0(\cal1_v__reg[7]|Q_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_abc_1582_), .F3(dummy_abc_1583_) );
      defparam ii2677.CONFIG_DATA = 16'h6666;
      defparam ii2677.PLACE_LOCATION = "NONE";
      defparam ii2677.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2678 ( .DX(nn2678), .F0(\cal1_v__reg[8]|Q_net ), .F1(dummy_abc_1584_), .F2(dummy_abc_1585_), .F3(dummy_abc_1586_) );
      defparam ii2678.CONFIG_DATA = 16'hAAAA;
      defparam ii2678.PLACE_LOCATION = "NONE";
      defparam ii2678.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2679 ( .DX(nn2679), .F0(\cal1_v__reg[9]|Q_net ), .F1(dummy_abc_1587_), .F2(dummy_abc_1588_), .F3(dummy_abc_1589_) );
      defparam ii2679.CONFIG_DATA = 16'hAAAA;
      defparam ii2679.PLACE_LOCATION = "NONE";
      defparam ii2679.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2680 ( .DX(nn2680), .F0(\cal1_v__reg[10]|Q_net ), .F1(dummy_abc_1590_), .F2(dummy_abc_1591_), .F3(dummy_abc_1592_) );
      defparam ii2680.CONFIG_DATA = 16'hAAAA;
      defparam ii2680.PLACE_LOCATION = "NONE";
      defparam ii2680.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2681 ( .DX(nn2681), .F0(\cal1_v__reg[11]|Q_net ), .F1(dummy_abc_1593_), .F2(dummy_abc_1594_), .F3(dummy_abc_1595_) );
      defparam ii2681.CONFIG_DATA = 16'hAAAA;
      defparam ii2681.PLACE_LOCATION = "NONE";
      defparam ii2681.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2682 ( .DX(nn2682), .F0(\cal1_v__reg[12]|Q_net ), .F1(dummy_abc_1596_), .F2(dummy_abc_1597_), .F3(dummy_abc_1598_) );
      defparam ii2682.CONFIG_DATA = 16'hAAAA;
      defparam ii2682.PLACE_LOCATION = "NONE";
      defparam ii2682.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2683 ( .DX(nn2683), .F0(\cal1_v__reg[13]|Q_net ), .F1(dummy_abc_1599_), .F2(dummy_abc_1600_), .F3(dummy_abc_1601_) );
      defparam ii2683.CONFIG_DATA = 16'hAAAA;
      defparam ii2683.PLACE_LOCATION = "NONE";
      defparam ii2683.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2684 ( .DX(nn2684), .F0(\cal1_v__reg[14]|Q_net ), .F1(dummy_abc_1602_), .F2(dummy_abc_1603_), .F3(dummy_abc_1604_) );
      defparam ii2684.CONFIG_DATA = 16'hAAAA;
      defparam ii2684.PLACE_LOCATION = "NONE";
      defparam ii2684.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2685 ( .DX(nn2685), .F0(\cal1_v__reg[15]|Q_net ), .F1(dummy_abc_1605_), .F2(dummy_abc_1606_), .F3(dummy_abc_1607_) );
      defparam ii2685.CONFIG_DATA = 16'hAAAA;
      defparam ii2685.PLACE_LOCATION = "NONE";
      defparam ii2685.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2686 ( .DX(nn2686), .F0(\cal1_v__reg[16]|Q_net ), .F1(dummy_abc_1608_), .F2(dummy_abc_1609_), .F3(dummy_abc_1610_) );
      defparam ii2686.CONFIG_DATA = 16'hAAAA;
      defparam ii2686.PLACE_LOCATION = "NONE";
      defparam ii2686.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_0_ ( 
        .CA( {\cal1_v__reg[16]|Q_net , \cal1_v__reg[15]|Q_net , 
              \cal1_v__reg[14]|Q_net , \cal1_v__reg[13]|Q_net , \cal1_v__reg[12]|Q_net , 
              \cal1_v__reg[11]|Q_net , \cal1_v__reg[10]|Q_net , \cal1_v__reg[9]|Q_net , 
              \cal1_v__reg[8]|Q_net , \cal1_v__reg[7]|Q_net , \cal1_v__reg[6]|Q_net , 
              \cal1_v__reg[5]|Q_net , \cal1_v__reg[4]|Q_net , \cal1_v__reg[3]|Q_net , 
              \cal1_v__reg[2]|Q_net , \cal1_v__reg[1]|Q_net , \cal1_v__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_139_ ), 
        .DX( {nn2686, nn2685, nn2684, nn2683, nn2682, nn2681, nn2680, nn2679, 
              nn2678, nn2677, nn2676, nn2675, nn2674, nn2673, nn2672, nn2671, 
              nn2645} ), 
        .SUM( {\cal1_u128_XORCI_16|SUM_net , \cal1_u128_XORCI_15|SUM_net , 
              \cal1_u128_XORCI_14|SUM_net , \cal1_u128_XORCI_13|SUM_net , \cal1_u128_XORCI_12|SUM_net , 
              \cal1_u128_XORCI_11|SUM_net , \cal1_u128_XORCI_10|SUM_net , \cal1_u128_XORCI_9|SUM_net , 
              \cal1_u128_XORCI_8|SUM_net , \cal1_u128_XORCI_7|SUM_net , \cal1_u128_XORCI_6|SUM_net , 
              \cal1_u128_XORCI_5|SUM_net , \cal1_u128_XORCI_4|SUM_net , \cal1_u128_XORCI_3|SUM_net , 
              \cal1_u128_XORCI_2|SUM_net , \cal1_u128_XORCI_1|SUM_net , \cal1_u128_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2706 ( .DX(nn2706), .F0(\cal1_v__reg[6]|Q_net ), .F1(\cal1_u128_XORCI_6|SUM_net ), .F2(dummy_abc_1611_), .F3(dummy_abc_1612_) );
      defparam ii2706.CONFIG_DATA = 16'h2222;
      defparam ii2706.PLACE_LOCATION = "NONE";
      defparam ii2706.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2707 ( .DX(nn2707), .F0(\cal1_v__reg[8]|Q_net ), .F1(\cal1_u128_XORCI_8|SUM_net ), .F2(dummy_abc_1613_), .F3(dummy_abc_1614_) );
      defparam ii2707.CONFIG_DATA = 16'h6666;
      defparam ii2707.PLACE_LOCATION = "NONE";
      defparam ii2707.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2708 ( .DX(nn2708), .F0(\cal1_v__reg[7]|Q_net ), .F1(\cal1_u128_XORCI_7|SUM_net ), .F2(nn2706), .F3(nn2707) );
      defparam ii2708.CONFIG_DATA = 16'hDFB6;
      defparam ii2708.PLACE_LOCATION = "NONE";
      defparam ii2708.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2709 ( .DX(nn2709), .F0(\cal1_v__reg[6]|Q_net ), .F1(dummy_123_), .F2(\cal1_u128_XORCI_6|SUM_net ), .F3(nn1328) );
      defparam ii2709.CONFIG_DATA = 16'h1200;
      defparam ii2709.PLACE_LOCATION = "NONE";
      defparam ii2709.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2710 ( .DX(nn2710), .F0(dummy_35_), .F1(nn1331), .F2(nn2708), .F3(nn2709) );
      defparam ii2710.CONFIG_DATA = 16'h1F11;
      defparam ii2710.PLACE_LOCATION = "NONE";
      defparam ii2710.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2711 ( .DX(nn2711), .F0(dummy_123_), .F1(dummy_35_), .F2(dummy_22_), .F3(nn2708) );
      defparam ii2711.CONFIG_DATA = 16'h0400;
      defparam ii2711.PLACE_LOCATION = "NONE";
      defparam ii2711.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2712 ( .DX(nn2712), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1615_), .F3(dummy_abc_1616_) );
      defparam ii2712.CONFIG_DATA = 16'h9999;
      defparam ii2712.PLACE_LOCATION = "NONE";
      defparam ii2712.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2713 ( .DX(nn2713), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1617_), .F3(dummy_abc_1618_) );
      defparam ii2713.CONFIG_DATA = 16'h9999;
      defparam ii2713.PLACE_LOCATION = "NONE";
      defparam ii2713.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2714 ( .DX(nn2714), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_abc_1619_), .F3(dummy_abc_1620_) );
      defparam ii2714.CONFIG_DATA = 16'h9999;
      defparam ii2714.PLACE_LOCATION = "NONE";
      defparam ii2714.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2715 ( .DX(nn2715), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[3]|Q_net ), .F2(dummy_abc_1621_), .F3(dummy_abc_1622_) );
      defparam ii2715.CONFIG_DATA = 16'h9999;
      defparam ii2715.PLACE_LOCATION = "NONE";
      defparam ii2715.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2716 ( .DX(nn2716), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[4]|Q_net ), .F2(dummy_abc_1623_), .F3(dummy_abc_1624_) );
      defparam ii2716.CONFIG_DATA = 16'h9999;
      defparam ii2716.PLACE_LOCATION = "NONE";
      defparam ii2716.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2717 ( .DX(nn2717), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[5]|Q_net ), .F2(dummy_abc_1625_), .F3(dummy_abc_1626_) );
      defparam ii2717.CONFIG_DATA = 16'h9999;
      defparam ii2717.PLACE_LOCATION = "NONE";
      defparam ii2717.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2718 ( .DX(nn2718), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[6]|Q_net ), .F2(dummy_abc_1627_), .F3(dummy_abc_1628_) );
      defparam ii2718.CONFIG_DATA = 16'h9999;
      defparam ii2718.PLACE_LOCATION = "NONE";
      defparam ii2718.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2719 ( .DX(nn2719), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[7]|Q_net ), .F2(dummy_abc_1629_), .F3(dummy_abc_1630_) );
      defparam ii2719.CONFIG_DATA = 16'h9999;
      defparam ii2719.PLACE_LOCATION = "NONE";
      defparam ii2719.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2720 ( .DX(nn2720), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[8]|Q_net ), .F2(dummy_abc_1631_), .F3(dummy_abc_1632_) );
      defparam ii2720.CONFIG_DATA = 16'h9999;
      defparam ii2720.PLACE_LOCATION = "NONE";
      defparam ii2720.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2721 ( .DX(nn2721), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[9]|Q_net ), .F2(dummy_abc_1633_), .F3(dummy_abc_1634_) );
      defparam ii2721.CONFIG_DATA = 16'h9999;
      defparam ii2721.PLACE_LOCATION = "NONE";
      defparam ii2721.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2722 ( .DX(nn2722), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[10]|Q_net ), .F2(dummy_abc_1635_), .F3(dummy_abc_1636_) );
      defparam ii2722.CONFIG_DATA = 16'h9999;
      defparam ii2722.PLACE_LOCATION = "NONE";
      defparam ii2722.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2723 ( .DX(nn2723), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[11]|Q_net ), .F2(dummy_abc_1637_), .F3(dummy_abc_1638_) );
      defparam ii2723.CONFIG_DATA = 16'h9999;
      defparam ii2723.PLACE_LOCATION = "NONE";
      defparam ii2723.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2724 ( .DX(nn2724), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[12]|Q_net ), .F2(dummy_abc_1639_), .F3(dummy_abc_1640_) );
      defparam ii2724.CONFIG_DATA = 16'h9999;
      defparam ii2724.PLACE_LOCATION = "NONE";
      defparam ii2724.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2725 ( .DX(nn2725), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[13]|Q_net ), .F2(dummy_abc_1641_), .F3(dummy_abc_1642_) );
      defparam ii2725.CONFIG_DATA = 16'h9999;
      defparam ii2725.PLACE_LOCATION = "NONE";
      defparam ii2725.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2726 ( .DX(nn2726), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[14]|Q_net ), .F2(dummy_abc_1643_), .F3(dummy_abc_1644_) );
      defparam ii2726.CONFIG_DATA = 16'h9999;
      defparam ii2726.PLACE_LOCATION = "NONE";
      defparam ii2726.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2727 ( .DX(nn2727), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[15]|Q_net ), .F2(dummy_abc_1645_), .F3(dummy_abc_1646_) );
      defparam ii2727.CONFIG_DATA = 16'h9999;
      defparam ii2727.PLACE_LOCATION = "NONE";
      defparam ii2727.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2728 ( .DX(nn2728), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1647_), .F3(dummy_abc_1648_) );
      defparam ii2728.CONFIG_DATA = 16'h9999;
      defparam ii2728.PLACE_LOCATION = "NONE";
      defparam ii2728.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2729 ( .DX(nn2729), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1649_), .F3(dummy_abc_1650_) );
      defparam ii2729.CONFIG_DATA = 16'h9999;
      defparam ii2729.PLACE_LOCATION = "NONE";
      defparam ii2729.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2730 ( .DX(nn2730), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1651_), .F3(dummy_abc_1652_) );
      defparam ii2730.CONFIG_DATA = 16'h9999;
      defparam ii2730.PLACE_LOCATION = "NONE";
      defparam ii2730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2731 ( .DX(nn2731), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_abc_1653_), .F2(dummy_abc_1654_), .F3(dummy_abc_1655_) );
      defparam ii2731.CONFIG_DATA = 16'h5555;
      defparam ii2731.PLACE_LOCATION = "NONE";
      defparam ii2731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2732 ( .DX(nn2732), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1656_), .F2(dummy_abc_1657_), .F3(dummy_abc_1658_) );
      defparam ii2732.CONFIG_DATA = 16'h5555;
      defparam ii2732.PLACE_LOCATION = "NONE";
      defparam ii2732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2733 ( .DX(nn2733), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1659_), .F2(dummy_abc_1660_), .F3(dummy_abc_1661_) );
      defparam ii2733.CONFIG_DATA = 16'h5555;
      defparam ii2733.PLACE_LOCATION = "NONE";
      defparam ii2733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2734 ( .DX(nn2734), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1662_), .F2(dummy_abc_1663_), .F3(dummy_abc_1664_) );
      defparam ii2734.CONFIG_DATA = 16'h5555;
      defparam ii2734.PLACE_LOCATION = "NONE";
      defparam ii2734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2735 ( .DX(nn2735), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1665_), .F2(dummy_abc_1666_), .F3(dummy_abc_1667_) );
      defparam ii2735.CONFIG_DATA = 16'h5555;
      defparam ii2735.PLACE_LOCATION = "NONE";
      defparam ii2735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2736 ( .DX(nn2736), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1668_), .F2(dummy_abc_1669_), .F3(dummy_abc_1670_) );
      defparam ii2736.CONFIG_DATA = 16'h5555;
      defparam ii2736.PLACE_LOCATION = "NONE";
      defparam ii2736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2737 ( .DX(nn2737), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1671_), .F2(dummy_abc_1672_), .F3(dummy_abc_1673_) );
      defparam ii2737.CONFIG_DATA = 16'h5555;
      defparam ii2737.PLACE_LOCATION = "NONE";
      defparam ii2737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2738 ( .DX(nn2738), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1674_), .F2(dummy_abc_1675_), .F3(dummy_abc_1676_) );
      defparam ii2738.CONFIG_DATA = 16'h5555;
      defparam ii2738.PLACE_LOCATION = "NONE";
      defparam ii2738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2739 ( .DX(nn2739), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1677_), .F2(dummy_abc_1678_), .F3(dummy_abc_1679_) );
      defparam ii2739.CONFIG_DATA = 16'h5555;
      defparam ii2739.PLACE_LOCATION = "NONE";
      defparam ii2739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2740 ( .DX(nn2740), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1680_), .F2(dummy_abc_1681_), .F3(dummy_abc_1682_) );
      defparam ii2740.CONFIG_DATA = 16'h5555;
      defparam ii2740.PLACE_LOCATION = "NONE";
      defparam ii2740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2741 ( .DX(nn2741), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1683_), .F2(dummy_abc_1684_), .F3(dummy_abc_1685_) );
      defparam ii2741.CONFIG_DATA = 16'h5555;
      defparam ii2741.PLACE_LOCATION = "NONE";
      defparam ii2741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2742 ( .DX(nn2742), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1686_), .F2(dummy_abc_1687_), .F3(dummy_abc_1688_) );
      defparam ii2742.CONFIG_DATA = 16'h5555;
      defparam ii2742.PLACE_LOCATION = "NONE";
      defparam ii2742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2743 ( .DX(nn2743), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1689_), .F2(dummy_abc_1690_), .F3(dummy_abc_1691_) );
      defparam ii2743.CONFIG_DATA = 16'h5555;
      defparam ii2743.PLACE_LOCATION = "NONE";
      defparam ii2743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2744 ( .DX(nn2744), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1692_), .F2(dummy_abc_1693_), .F3(dummy_abc_1694_) );
      defparam ii2744.CONFIG_DATA = 16'h5555;
      defparam ii2744.PLACE_LOCATION = "NONE";
      defparam ii2744.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2745 ( .DX(nn2745), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1695_), .F2(dummy_abc_1696_), .F3(dummy_abc_1697_) );
      defparam ii2745.CONFIG_DATA = 16'h5555;
      defparam ii2745.PLACE_LOCATION = "NONE";
      defparam ii2745.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2746 ( .DX(nn2746), .F0(dummy_abc_1698_), .F1(dummy_abc_1699_), .F2(dummy_abc_1700_), .F3(dummy_abc_1701_) );
      defparam ii2746.CONFIG_DATA = 16'hFFFF;
      defparam ii2746.PLACE_LOCATION = "NONE";
      defparam ii2746.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_24_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_222_ ), 
        .DX( {nn2746, nn2745, nn2744, nn2743, nn2742, nn2741, nn2740, nn2739, 
              nn2738, nn2737, nn2736, nn2735, nn2734, nn2733, nn2732, nn2731, 
              nn2730, nn2729} ), 
        .SUM( {\coefcal1_divide_inst1_u120_XORCI_17|SUM_net , dummy_223_, 
              dummy_224_, dummy_225_, dummy_226_, dummy_227_, dummy_228_, dummy_229_, 
              dummy_230_, dummy_231_, dummy_232_, dummy_233_, dummy_234_, dummy_235_, 
              dummy_236_, dummy_237_, dummy_238_, dummy_239_} )
      );
    CS_LUT4_PRIM ii2767 ( .DX(nn2767), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_222_) );
      defparam ii2767.CONFIG_DATA = 16'hA569;
      defparam ii2767.PLACE_LOCATION = "NONE";
      defparam ii2767.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2768 ( .DX(nn2768), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1702_), .F3(dummy_abc_1703_) );
      defparam ii2768.CONFIG_DATA = 16'h9999;
      defparam ii2768.PLACE_LOCATION = "NONE";
      defparam ii2768.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2769 ( .DX(nn2769), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1704_), .F3(dummy_abc_1705_) );
      defparam ii2769.CONFIG_DATA = 16'h9999;
      defparam ii2769.PLACE_LOCATION = "NONE";
      defparam ii2769.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2770 ( .DX(nn2770), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_abc_1706_), .F2(dummy_abc_1707_), .F3(dummy_abc_1708_) );
      defparam ii2770.CONFIG_DATA = 16'h5555;
      defparam ii2770.PLACE_LOCATION = "NONE";
      defparam ii2770.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2771 ( .DX(nn2771), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1709_), .F2(dummy_abc_1710_), .F3(dummy_abc_1711_) );
      defparam ii2771.CONFIG_DATA = 16'h5555;
      defparam ii2771.PLACE_LOCATION = "NONE";
      defparam ii2771.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2772 ( .DX(nn2772), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1712_), .F2(dummy_abc_1713_), .F3(dummy_abc_1714_) );
      defparam ii2772.CONFIG_DATA = 16'h5555;
      defparam ii2772.PLACE_LOCATION = "NONE";
      defparam ii2772.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2773 ( .DX(nn2773), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1715_), .F2(dummy_abc_1716_), .F3(dummy_abc_1717_) );
      defparam ii2773.CONFIG_DATA = 16'h5555;
      defparam ii2773.PLACE_LOCATION = "NONE";
      defparam ii2773.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2774 ( .DX(nn2774), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1718_), .F2(dummy_abc_1719_), .F3(dummy_abc_1720_) );
      defparam ii2774.CONFIG_DATA = 16'h5555;
      defparam ii2774.PLACE_LOCATION = "NONE";
      defparam ii2774.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2775 ( .DX(nn2775), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1721_), .F2(dummy_abc_1722_), .F3(dummy_abc_1723_) );
      defparam ii2775.CONFIG_DATA = 16'h5555;
      defparam ii2775.PLACE_LOCATION = "NONE";
      defparam ii2775.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2776 ( .DX(nn2776), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1724_), .F2(dummy_abc_1725_), .F3(dummy_abc_1726_) );
      defparam ii2776.CONFIG_DATA = 16'h5555;
      defparam ii2776.PLACE_LOCATION = "NONE";
      defparam ii2776.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2777 ( .DX(nn2777), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1727_), .F2(dummy_abc_1728_), .F3(dummy_abc_1729_) );
      defparam ii2777.CONFIG_DATA = 16'h5555;
      defparam ii2777.PLACE_LOCATION = "NONE";
      defparam ii2777.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2778 ( .DX(nn2778), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1730_), .F2(dummy_abc_1731_), .F3(dummy_abc_1732_) );
      defparam ii2778.CONFIG_DATA = 16'h5555;
      defparam ii2778.PLACE_LOCATION = "NONE";
      defparam ii2778.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2779 ( .DX(nn2779), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1733_), .F2(dummy_abc_1734_), .F3(dummy_abc_1735_) );
      defparam ii2779.CONFIG_DATA = 16'h5555;
      defparam ii2779.PLACE_LOCATION = "NONE";
      defparam ii2779.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2780 ( .DX(nn2780), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1736_), .F2(dummy_abc_1737_), .F3(dummy_abc_1738_) );
      defparam ii2780.CONFIG_DATA = 16'h5555;
      defparam ii2780.PLACE_LOCATION = "NONE";
      defparam ii2780.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2781 ( .DX(nn2781), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1739_), .F2(dummy_abc_1740_), .F3(dummy_abc_1741_) );
      defparam ii2781.CONFIG_DATA = 16'h5555;
      defparam ii2781.PLACE_LOCATION = "NONE";
      defparam ii2781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2782 ( .DX(nn2782), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1742_), .F2(dummy_abc_1743_), .F3(dummy_abc_1744_) );
      defparam ii2782.CONFIG_DATA = 16'h5555;
      defparam ii2782.PLACE_LOCATION = "NONE";
      defparam ii2782.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2783 ( .DX(nn2783), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1745_), .F2(dummy_abc_1746_), .F3(dummy_abc_1747_) );
      defparam ii2783.CONFIG_DATA = 16'h5555;
      defparam ii2783.PLACE_LOCATION = "NONE";
      defparam ii2783.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2784 ( .DX(nn2784), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1748_), .F2(dummy_abc_1749_), .F3(dummy_abc_1750_) );
      defparam ii2784.CONFIG_DATA = 16'h5555;
      defparam ii2784.PLACE_LOCATION = "NONE";
      defparam ii2784.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_9_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, \coefcal1_xDividend__reg[16]|Q_net , 
              \coefcal1_xDividend__reg[15]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_200_ ), 
        .DX( {nn2784, nn2783, nn2782, nn2781, nn2780, nn2779, nn2778, nn2777, 
              nn2776, nn2775, nn2774, nn2773, nn2772, nn2771, nn2770, nn2769, 
              nn2768} ), 
        .SUM( {dummy_201_, \coefcal1_divide_inst1_u102_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_14|SUM_net , \coefcal1_divide_inst1_u102_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_12|SUM_net , \coefcal1_divide_inst1_u102_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_10|SUM_net , \coefcal1_divide_inst1_u102_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_8|SUM_net , \coefcal1_divide_inst1_u102_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_6|SUM_net , \coefcal1_divide_inst1_u102_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_4|SUM_net , \coefcal1_divide_inst1_u102_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_2|SUM_net , \coefcal1_divide_inst1_u102_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2804 ( .DX(nn2804), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_222_), .F3(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ) );
      defparam ii2804.CONFIG_DATA = 16'h9C93;
      defparam ii2804.PLACE_LOCATION = "NONE";
      defparam ii2804.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2805 ( .DX(nn2805), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1751_), .F2(dummy_abc_1752_), .F3(dummy_abc_1753_) );
      defparam ii2805.CONFIG_DATA = 16'h5555;
      defparam ii2805.PLACE_LOCATION = "NONE";
      defparam ii2805.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2806 ( .DX(nn2806), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1754_), .F2(dummy_abc_1755_), .F3(dummy_abc_1756_) );
      defparam ii2806.CONFIG_DATA = 16'h5555;
      defparam ii2806.PLACE_LOCATION = "NONE";
      defparam ii2806.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2807 ( .DX(nn2807), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1757_), .F2(dummy_abc_1758_), .F3(dummy_abc_1759_) );
      defparam ii2807.CONFIG_DATA = 16'h5555;
      defparam ii2807.PLACE_LOCATION = "NONE";
      defparam ii2807.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2808 ( .DX(nn2808), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1760_), .F2(dummy_abc_1761_), .F3(dummy_abc_1762_) );
      defparam ii2808.CONFIG_DATA = 16'h5555;
      defparam ii2808.PLACE_LOCATION = "NONE";
      defparam ii2808.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2809 ( .DX(nn2809), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1763_), .F2(dummy_abc_1764_), .F3(dummy_abc_1765_) );
      defparam ii2809.CONFIG_DATA = 16'h5555;
      defparam ii2809.PLACE_LOCATION = "NONE";
      defparam ii2809.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2810 ( .DX(nn2810), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1766_), .F2(dummy_abc_1767_), .F3(dummy_abc_1768_) );
      defparam ii2810.CONFIG_DATA = 16'h5555;
      defparam ii2810.PLACE_LOCATION = "NONE";
      defparam ii2810.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2811 ( .DX(nn2811), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1769_), .F2(dummy_abc_1770_), .F3(dummy_abc_1771_) );
      defparam ii2811.CONFIG_DATA = 16'h5555;
      defparam ii2811.PLACE_LOCATION = "NONE";
      defparam ii2811.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2812 ( .DX(nn2812), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1772_), .F2(dummy_abc_1773_), .F3(dummy_abc_1774_) );
      defparam ii2812.CONFIG_DATA = 16'h5555;
      defparam ii2812.PLACE_LOCATION = "NONE";
      defparam ii2812.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2813 ( .DX(nn2813), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1775_), .F2(dummy_abc_1776_), .F3(dummy_abc_1777_) );
      defparam ii2813.CONFIG_DATA = 16'h5555;
      defparam ii2813.PLACE_LOCATION = "NONE";
      defparam ii2813.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2814 ( .DX(nn2814), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1778_), .F2(dummy_abc_1779_), .F3(dummy_abc_1780_) );
      defparam ii2814.CONFIG_DATA = 16'h5555;
      defparam ii2814.PLACE_LOCATION = "NONE";
      defparam ii2814.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2815 ( .DX(nn2815), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1781_), .F2(dummy_abc_1782_), .F3(dummy_abc_1783_) );
      defparam ii2815.CONFIG_DATA = 16'h5555;
      defparam ii2815.PLACE_LOCATION = "NONE";
      defparam ii2815.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2816 ( .DX(nn2816), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1784_), .F2(dummy_abc_1785_), .F3(dummy_abc_1786_) );
      defparam ii2816.CONFIG_DATA = 16'h5555;
      defparam ii2816.PLACE_LOCATION = "NONE";
      defparam ii2816.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2817 ( .DX(nn2817), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1787_), .F2(dummy_abc_1788_), .F3(dummy_abc_1789_) );
      defparam ii2817.CONFIG_DATA = 16'h5555;
      defparam ii2817.PLACE_LOCATION = "NONE";
      defparam ii2817.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2818 ( .DX(nn2818), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1790_), .F2(dummy_abc_1791_), .F3(dummy_abc_1792_) );
      defparam ii2818.CONFIG_DATA = 16'h5555;
      defparam ii2818.PLACE_LOCATION = "NONE";
      defparam ii2818.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2819 ( .DX(nn2819), .F0(dummy_abc_1793_), .F1(dummy_abc_1794_), .F2(dummy_abc_1795_), .F3(dummy_abc_1796_) );
      defparam ii2819.CONFIG_DATA = 16'hFFFF;
      defparam ii2819.PLACE_LOCATION = "NONE";
      defparam ii2819.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_25_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_241_ ), 
        .DX( {nn2819, nn2818, nn2817, nn2816, nn2815, nn2814, nn2813, nn2812, 
              nn2811, nn2810, nn2809, nn2808, nn2807, nn2806, nn2805, nn2804, 
              nn2767, nn2728} ), 
        .SUM( {\coefcal1_divide_inst1_u122_XORCI_17|SUM_net , dummy_242_, 
              dummy_243_, dummy_244_, dummy_245_, dummy_246_, dummy_247_, dummy_248_, 
              dummy_249_, dummy_250_, dummy_251_, dummy_252_, dummy_253_, dummy_254_, 
              dummy_255_, dummy_256_, dummy_257_, dummy_258_} )
      );
    CS_LUT4_PRIM ii2840 ( .DX(nn2840), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1797_), .F3(dummy_abc_1798_) );
      defparam ii2840.CONFIG_DATA = 16'h9999;
      defparam ii2840.PLACE_LOCATION = "NONE";
      defparam ii2840.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2841 ( .DX(nn2841), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_241_) );
      defparam ii2841.CONFIG_DATA = 16'hA569;
      defparam ii2841.PLACE_LOCATION = "NONE";
      defparam ii2841.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2842 ( .DX(nn2842), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_222_), .F3(dummy_abc_1799_) );
      defparam ii2842.CONFIG_DATA = 16'hA6A6;
      defparam ii2842.PLACE_LOCATION = "NONE";
      defparam ii2842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2843 ( .DX(nn2843), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(dummy_222_), .F2(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ), .F3(dummy_abc_1800_) );
      defparam ii2843.CONFIG_DATA = 16'hB8B8;
      defparam ii2843.PLACE_LOCATION = "NONE";
      defparam ii2843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2844 ( .DX(nn2844), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1801_), .F3(dummy_abc_1802_) );
      defparam ii2844.CONFIG_DATA = 16'h9999;
      defparam ii2844.PLACE_LOCATION = "NONE";
      defparam ii2844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2845 ( .DX(nn2845), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_222_) );
      defparam ii2845.CONFIG_DATA = 16'hA569;
      defparam ii2845.PLACE_LOCATION = "NONE";
      defparam ii2845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2846 ( .DX(nn2846), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_222_), .F3(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ) );
      defparam ii2846.CONFIG_DATA = 16'h9C93;
      defparam ii2846.PLACE_LOCATION = "NONE";
      defparam ii2846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2847 ( .DX(nn2847), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1803_), .F2(dummy_abc_1804_), .F3(dummy_abc_1805_) );
      defparam ii2847.CONFIG_DATA = 16'h5555;
      defparam ii2847.PLACE_LOCATION = "NONE";
      defparam ii2847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2848 ( .DX(nn2848), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1806_), .F2(dummy_abc_1807_), .F3(dummy_abc_1808_) );
      defparam ii2848.CONFIG_DATA = 16'h5555;
      defparam ii2848.PLACE_LOCATION = "NONE";
      defparam ii2848.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2849 ( .DX(nn2849), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1809_), .F2(dummy_abc_1810_), .F3(dummy_abc_1811_) );
      defparam ii2849.CONFIG_DATA = 16'h5555;
      defparam ii2849.PLACE_LOCATION = "NONE";
      defparam ii2849.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2850 ( .DX(nn2850), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1812_), .F2(dummy_abc_1813_), .F3(dummy_abc_1814_) );
      defparam ii2850.CONFIG_DATA = 16'h5555;
      defparam ii2850.PLACE_LOCATION = "NONE";
      defparam ii2850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2851 ( .DX(nn2851), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1815_), .F2(dummy_abc_1816_), .F3(dummy_abc_1817_) );
      defparam ii2851.CONFIG_DATA = 16'h5555;
      defparam ii2851.PLACE_LOCATION = "NONE";
      defparam ii2851.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2852 ( .DX(nn2852), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1818_), .F2(dummy_abc_1819_), .F3(dummy_abc_1820_) );
      defparam ii2852.CONFIG_DATA = 16'h5555;
      defparam ii2852.PLACE_LOCATION = "NONE";
      defparam ii2852.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2853 ( .DX(nn2853), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1821_), .F2(dummy_abc_1822_), .F3(dummy_abc_1823_) );
      defparam ii2853.CONFIG_DATA = 16'h5555;
      defparam ii2853.PLACE_LOCATION = "NONE";
      defparam ii2853.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2854 ( .DX(nn2854), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1824_), .F2(dummy_abc_1825_), .F3(dummy_abc_1826_) );
      defparam ii2854.CONFIG_DATA = 16'h5555;
      defparam ii2854.PLACE_LOCATION = "NONE";
      defparam ii2854.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2855 ( .DX(nn2855), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1827_), .F2(dummy_abc_1828_), .F3(dummy_abc_1829_) );
      defparam ii2855.CONFIG_DATA = 16'h5555;
      defparam ii2855.PLACE_LOCATION = "NONE";
      defparam ii2855.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2856 ( .DX(nn2856), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1830_), .F2(dummy_abc_1831_), .F3(dummy_abc_1832_) );
      defparam ii2856.CONFIG_DATA = 16'h5555;
      defparam ii2856.PLACE_LOCATION = "NONE";
      defparam ii2856.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2857 ( .DX(nn2857), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1833_), .F2(dummy_abc_1834_), .F3(dummy_abc_1835_) );
      defparam ii2857.CONFIG_DATA = 16'h5555;
      defparam ii2857.PLACE_LOCATION = "NONE";
      defparam ii2857.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2858 ( .DX(nn2858), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1836_), .F2(dummy_abc_1837_), .F3(dummy_abc_1838_) );
      defparam ii2858.CONFIG_DATA = 16'h5555;
      defparam ii2858.PLACE_LOCATION = "NONE";
      defparam ii2858.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2859 ( .DX(nn2859), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1839_), .F2(dummy_abc_1840_), .F3(dummy_abc_1841_) );
      defparam ii2859.CONFIG_DATA = 16'h5555;
      defparam ii2859.PLACE_LOCATION = "NONE";
      defparam ii2859.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2860 ( .DX(nn2860), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1842_), .F2(dummy_abc_1843_), .F3(dummy_abc_1844_) );
      defparam ii2860.CONFIG_DATA = 16'h5555;
      defparam ii2860.PLACE_LOCATION = "NONE";
      defparam ii2860.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_10_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2843, 
              nn2842, \coefcal1_xDividend__reg[14]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_140_ ), 
        .DX( {nn2860, nn2859, nn2858, nn2857, nn2856, nn2855, nn2854, nn2853, 
              nn2852, nn2851, nn2850, nn2849, nn2848, nn2847, nn2846, nn2845, 
              nn2844} ), 
        .SUM( {dummy_141_, \coefcal1_divide_inst1_u103_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_14|SUM_net , \coefcal1_divide_inst1_u103_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_12|SUM_net , \coefcal1_divide_inst1_u103_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_10|SUM_net , \coefcal1_divide_inst1_u103_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_8|SUM_net , \coefcal1_divide_inst1_u103_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_6|SUM_net , \coefcal1_divide_inst1_u103_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_4|SUM_net , \coefcal1_divide_inst1_u103_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_2|SUM_net , \coefcal1_divide_inst1_u103_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2880 ( .DX(nn2880), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_241_), .F2(nn2842), .F3(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ) );
      defparam ii2880.CONFIG_DATA = 16'hA695;
      defparam ii2880.PLACE_LOCATION = "NONE";
      defparam ii2880.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2881 ( .DX(nn2881), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2843), .F2(dummy_241_), .F3(\coefcal1_divide_inst1_u103_XORCI_2|SUM_net ) );
      defparam ii2881.CONFIG_DATA = 16'h9A95;
      defparam ii2881.PLACE_LOCATION = "NONE";
      defparam ii2881.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2882 ( .DX(nn2882), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1845_), .F2(dummy_abc_1846_), .F3(dummy_abc_1847_) );
      defparam ii2882.CONFIG_DATA = 16'h5555;
      defparam ii2882.PLACE_LOCATION = "NONE";
      defparam ii2882.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2883 ( .DX(nn2883), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1848_), .F2(dummy_abc_1849_), .F3(dummy_abc_1850_) );
      defparam ii2883.CONFIG_DATA = 16'h5555;
      defparam ii2883.PLACE_LOCATION = "NONE";
      defparam ii2883.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2884 ( .DX(nn2884), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1851_), .F2(dummy_abc_1852_), .F3(dummy_abc_1853_) );
      defparam ii2884.CONFIG_DATA = 16'h5555;
      defparam ii2884.PLACE_LOCATION = "NONE";
      defparam ii2884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2885 ( .DX(nn2885), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1854_), .F2(dummy_abc_1855_), .F3(dummy_abc_1856_) );
      defparam ii2885.CONFIG_DATA = 16'h5555;
      defparam ii2885.PLACE_LOCATION = "NONE";
      defparam ii2885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2886 ( .DX(nn2886), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1857_), .F2(dummy_abc_1858_), .F3(dummy_abc_1859_) );
      defparam ii2886.CONFIG_DATA = 16'h5555;
      defparam ii2886.PLACE_LOCATION = "NONE";
      defparam ii2886.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2887 ( .DX(nn2887), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1860_), .F2(dummy_abc_1861_), .F3(dummy_abc_1862_) );
      defparam ii2887.CONFIG_DATA = 16'h5555;
      defparam ii2887.PLACE_LOCATION = "NONE";
      defparam ii2887.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2888 ( .DX(nn2888), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1863_), .F2(dummy_abc_1864_), .F3(dummy_abc_1865_) );
      defparam ii2888.CONFIG_DATA = 16'h5555;
      defparam ii2888.PLACE_LOCATION = "NONE";
      defparam ii2888.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2889 ( .DX(nn2889), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1866_), .F2(dummy_abc_1867_), .F3(dummy_abc_1868_) );
      defparam ii2889.CONFIG_DATA = 16'h5555;
      defparam ii2889.PLACE_LOCATION = "NONE";
      defparam ii2889.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2890 ( .DX(nn2890), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1869_), .F2(dummy_abc_1870_), .F3(dummy_abc_1871_) );
      defparam ii2890.CONFIG_DATA = 16'h5555;
      defparam ii2890.PLACE_LOCATION = "NONE";
      defparam ii2890.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2891 ( .DX(nn2891), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1872_), .F2(dummy_abc_1873_), .F3(dummy_abc_1874_) );
      defparam ii2891.CONFIG_DATA = 16'h5555;
      defparam ii2891.PLACE_LOCATION = "NONE";
      defparam ii2891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2892 ( .DX(nn2892), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1875_), .F2(dummy_abc_1876_), .F3(dummy_abc_1877_) );
      defparam ii2892.CONFIG_DATA = 16'h5555;
      defparam ii2892.PLACE_LOCATION = "NONE";
      defparam ii2892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2893 ( .DX(nn2893), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1878_), .F2(dummy_abc_1879_), .F3(dummy_abc_1880_) );
      defparam ii2893.CONFIG_DATA = 16'h5555;
      defparam ii2893.PLACE_LOCATION = "NONE";
      defparam ii2893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2894 ( .DX(nn2894), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1881_), .F2(dummy_abc_1882_), .F3(dummy_abc_1883_) );
      defparam ii2894.CONFIG_DATA = 16'h5555;
      defparam ii2894.PLACE_LOCATION = "NONE";
      defparam ii2894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2895 ( .DX(nn2895), .F0(dummy_abc_1884_), .F1(dummy_abc_1885_), .F2(dummy_abc_1886_), .F3(dummy_abc_1887_) );
      defparam ii2895.CONFIG_DATA = 16'hFFFF;
      defparam ii2895.PLACE_LOCATION = "NONE";
      defparam ii2895.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_26_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_260_ ), 
        .DX( {nn2895, nn2894, nn2893, nn2892, nn2891, nn2890, nn2889, nn2888, 
              nn2887, nn2886, nn2885, nn2884, nn2883, nn2882, nn2881, nn2880, 
              nn2841, nn2840} ), 
        .SUM( {\coefcal1_divide_inst1_u124_XORCI_17|SUM_net , dummy_261_, 
              dummy_262_, dummy_263_, dummy_264_, dummy_265_, dummy_266_, dummy_267_, 
              dummy_268_, dummy_269_, dummy_270_, dummy_271_, dummy_272_, dummy_273_, 
              dummy_274_, dummy_275_, dummy_276_, dummy_277_} )
      );
    CS_LUT4_PRIM ii2916 ( .DX(nn2916), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_241_), .F3(dummy_abc_1888_) );
      defparam ii2916.CONFIG_DATA = 16'hA6A6;
      defparam ii2916.PLACE_LOCATION = "NONE";
      defparam ii2916.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2917 ( .DX(nn2917), .F0(dummy_241_), .F1(nn2842), .F2(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ), .F3(dummy_abc_1889_) );
      defparam ii2917.CONFIG_DATA = 16'hD8D8;
      defparam ii2917.PLACE_LOCATION = "NONE";
      defparam ii2917.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2918 ( .DX(nn2918), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1890_), .F3(dummy_abc_1891_) );
      defparam ii2918.CONFIG_DATA = 16'h9999;
      defparam ii2918.PLACE_LOCATION = "NONE";
      defparam ii2918.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2919 ( .DX(nn2919), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_241_) );
      defparam ii2919.CONFIG_DATA = 16'hA569;
      defparam ii2919.PLACE_LOCATION = "NONE";
      defparam ii2919.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2920 ( .DX(nn2920), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_241_), .F2(nn2842), .F3(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ) );
      defparam ii2920.CONFIG_DATA = 16'hA695;
      defparam ii2920.PLACE_LOCATION = "NONE";
      defparam ii2920.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2921 ( .DX(nn2921), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2843), .F2(dummy_241_), .F3(\coefcal1_divide_inst1_u103_XORCI_2|SUM_net ) );
      defparam ii2921.CONFIG_DATA = 16'h9A95;
      defparam ii2921.PLACE_LOCATION = "NONE";
      defparam ii2921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2922 ( .DX(nn2922), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1892_), .F2(dummy_abc_1893_), .F3(dummy_abc_1894_) );
      defparam ii2922.CONFIG_DATA = 16'h5555;
      defparam ii2922.PLACE_LOCATION = "NONE";
      defparam ii2922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2923 ( .DX(nn2923), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1895_), .F2(dummy_abc_1896_), .F3(dummy_abc_1897_) );
      defparam ii2923.CONFIG_DATA = 16'h5555;
      defparam ii2923.PLACE_LOCATION = "NONE";
      defparam ii2923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2924 ( .DX(nn2924), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1898_), .F2(dummy_abc_1899_), .F3(dummy_abc_1900_) );
      defparam ii2924.CONFIG_DATA = 16'h5555;
      defparam ii2924.PLACE_LOCATION = "NONE";
      defparam ii2924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2925 ( .DX(nn2925), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1901_), .F2(dummy_abc_1902_), .F3(dummy_abc_1903_) );
      defparam ii2925.CONFIG_DATA = 16'h5555;
      defparam ii2925.PLACE_LOCATION = "NONE";
      defparam ii2925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2926 ( .DX(nn2926), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1904_), .F2(dummy_abc_1905_), .F3(dummy_abc_1906_) );
      defparam ii2926.CONFIG_DATA = 16'h5555;
      defparam ii2926.PLACE_LOCATION = "NONE";
      defparam ii2926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2927 ( .DX(nn2927), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1907_), .F2(dummy_abc_1908_), .F3(dummy_abc_1909_) );
      defparam ii2927.CONFIG_DATA = 16'h5555;
      defparam ii2927.PLACE_LOCATION = "NONE";
      defparam ii2927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2928 ( .DX(nn2928), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1910_), .F2(dummy_abc_1911_), .F3(dummy_abc_1912_) );
      defparam ii2928.CONFIG_DATA = 16'h5555;
      defparam ii2928.PLACE_LOCATION = "NONE";
      defparam ii2928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2929 ( .DX(nn2929), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1913_), .F2(dummy_abc_1914_), .F3(dummy_abc_1915_) );
      defparam ii2929.CONFIG_DATA = 16'h5555;
      defparam ii2929.PLACE_LOCATION = "NONE";
      defparam ii2929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2930 ( .DX(nn2930), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1916_), .F2(dummy_abc_1917_), .F3(dummy_abc_1918_) );
      defparam ii2930.CONFIG_DATA = 16'h5555;
      defparam ii2930.PLACE_LOCATION = "NONE";
      defparam ii2930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2931 ( .DX(nn2931), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1919_), .F2(dummy_abc_1920_), .F3(dummy_abc_1921_) );
      defparam ii2931.CONFIG_DATA = 16'h5555;
      defparam ii2931.PLACE_LOCATION = "NONE";
      defparam ii2931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2932 ( .DX(nn2932), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1922_), .F2(dummy_abc_1923_), .F3(dummy_abc_1924_) );
      defparam ii2932.CONFIG_DATA = 16'h5555;
      defparam ii2932.PLACE_LOCATION = "NONE";
      defparam ii2932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2933 ( .DX(nn2933), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1925_), .F2(dummy_abc_1926_), .F3(dummy_abc_1927_) );
      defparam ii2933.CONFIG_DATA = 16'h5555;
      defparam ii2933.PLACE_LOCATION = "NONE";
      defparam ii2933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2934 ( .DX(nn2934), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1928_), .F2(dummy_abc_1929_), .F3(dummy_abc_1930_) );
      defparam ii2934.CONFIG_DATA = 16'h5555;
      defparam ii2934.PLACE_LOCATION = "NONE";
      defparam ii2934.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_11_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn2917, 
              nn2916, \coefcal1_xDividend__reg[13]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_142_ ), 
        .DX( {nn2934, nn2933, nn2932, nn2931, nn2930, nn2929, nn2928, nn2927, 
              nn2926, nn2925, nn2924, nn2923, nn2922, nn2921, nn2920, nn2919, 
              nn2918} ), 
        .SUM( {dummy_143_, \coefcal1_divide_inst1_u104_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_14|SUM_net , \coefcal1_divide_inst1_u104_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_12|SUM_net , \coefcal1_divide_inst1_u104_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_10|SUM_net , \coefcal1_divide_inst1_u104_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_8|SUM_net , \coefcal1_divide_inst1_u104_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_6|SUM_net , \coefcal1_divide_inst1_u104_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_4|SUM_net , \coefcal1_divide_inst1_u104_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_2|SUM_net , \coefcal1_divide_inst1_u104_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2954 ( .DX(nn2954), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(dummy_241_), .F2(dummy_260_), .F3(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ) );
      defparam ii2954.CONFIG_DATA = 16'h8F80;
      defparam ii2954.PLACE_LOCATION = "NONE";
      defparam ii2954.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2955 ( .DX(nn2955), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1931_), .F3(dummy_abc_1932_) );
      defparam ii2955.CONFIG_DATA = 16'h9999;
      defparam ii2955.PLACE_LOCATION = "NONE";
      defparam ii2955.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2956 ( .DX(nn2956), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_260_) );
      defparam ii2956.CONFIG_DATA = 16'hA569;
      defparam ii2956.PLACE_LOCATION = "NONE";
      defparam ii2956.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2957 ( .DX(nn2957), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_260_), .F2(nn2916), .F3(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ) );
      defparam ii2957.CONFIG_DATA = 16'hA695;
      defparam ii2957.PLACE_LOCATION = "NONE";
      defparam ii2957.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2958 ( .DX(nn2958), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2917), .F2(dummy_260_), .F3(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ) );
      defparam ii2958.CONFIG_DATA = 16'h9A95;
      defparam ii2958.PLACE_LOCATION = "NONE";
      defparam ii2958.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2959 ( .DX(nn2959), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[4]|Q_net ), .F2(dummy_241_), .F3(dummy_abc_1933_) );
      defparam ii2959.CONFIG_DATA = 16'h9393;
      defparam ii2959.PLACE_LOCATION = "NONE";
      defparam ii2959.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2960 ( .DX(nn2960), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_260_), .F2(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ), .F3(nn2959) );
      defparam ii2960.CONFIG_DATA = 16'hED21;
      defparam ii2960.PLACE_LOCATION = "NONE";
      defparam ii2960.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2961 ( .DX(nn2961), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1934_), .F2(dummy_abc_1935_), .F3(dummy_abc_1936_) );
      defparam ii2961.CONFIG_DATA = 16'h5555;
      defparam ii2961.PLACE_LOCATION = "NONE";
      defparam ii2961.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2962 ( .DX(nn2962), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1937_), .F2(dummy_abc_1938_), .F3(dummy_abc_1939_) );
      defparam ii2962.CONFIG_DATA = 16'h5555;
      defparam ii2962.PLACE_LOCATION = "NONE";
      defparam ii2962.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2963 ( .DX(nn2963), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1940_), .F2(dummy_abc_1941_), .F3(dummy_abc_1942_) );
      defparam ii2963.CONFIG_DATA = 16'h5555;
      defparam ii2963.PLACE_LOCATION = "NONE";
      defparam ii2963.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2964 ( .DX(nn2964), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1943_), .F2(dummy_abc_1944_), .F3(dummy_abc_1945_) );
      defparam ii2964.CONFIG_DATA = 16'h5555;
      defparam ii2964.PLACE_LOCATION = "NONE";
      defparam ii2964.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2965 ( .DX(nn2965), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1946_), .F2(dummy_abc_1947_), .F3(dummy_abc_1948_) );
      defparam ii2965.CONFIG_DATA = 16'h5555;
      defparam ii2965.PLACE_LOCATION = "NONE";
      defparam ii2965.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2966 ( .DX(nn2966), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1949_), .F2(dummy_abc_1950_), .F3(dummy_abc_1951_) );
      defparam ii2966.CONFIG_DATA = 16'h5555;
      defparam ii2966.PLACE_LOCATION = "NONE";
      defparam ii2966.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2967 ( .DX(nn2967), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1952_), .F2(dummy_abc_1953_), .F3(dummy_abc_1954_) );
      defparam ii2967.CONFIG_DATA = 16'h5555;
      defparam ii2967.PLACE_LOCATION = "NONE";
      defparam ii2967.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2968 ( .DX(nn2968), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1955_), .F2(dummy_abc_1956_), .F3(dummy_abc_1957_) );
      defparam ii2968.CONFIG_DATA = 16'h5555;
      defparam ii2968.PLACE_LOCATION = "NONE";
      defparam ii2968.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2969 ( .DX(nn2969), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1958_), .F2(dummy_abc_1959_), .F3(dummy_abc_1960_) );
      defparam ii2969.CONFIG_DATA = 16'h5555;
      defparam ii2969.PLACE_LOCATION = "NONE";
      defparam ii2969.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2970 ( .DX(nn2970), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1961_), .F2(dummy_abc_1962_), .F3(dummy_abc_1963_) );
      defparam ii2970.CONFIG_DATA = 16'h5555;
      defparam ii2970.PLACE_LOCATION = "NONE";
      defparam ii2970.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2971 ( .DX(nn2971), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1964_), .F2(dummy_abc_1965_), .F3(dummy_abc_1966_) );
      defparam ii2971.CONFIG_DATA = 16'h5555;
      defparam ii2971.PLACE_LOCATION = "NONE";
      defparam ii2971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2972 ( .DX(nn2972), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1967_), .F2(dummy_abc_1968_), .F3(dummy_abc_1969_) );
      defparam ii2972.CONFIG_DATA = 16'h5555;
      defparam ii2972.PLACE_LOCATION = "NONE";
      defparam ii2972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2973 ( .DX(nn2973), .F0(dummy_abc_1970_), .F1(dummy_abc_1971_), .F2(dummy_abc_1972_), .F3(dummy_abc_1973_) );
      defparam ii2973.CONFIG_DATA = 16'hFFFF;
      defparam ii2973.PLACE_LOCATION = "NONE";
      defparam ii2973.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_27_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_279_ ), 
        .DX( {nn2973, nn2972, nn2971, nn2970, nn2969, nn2968, nn2967, nn2966, 
              nn2965, nn2964, nn2963, nn2962, nn2961, nn2960, nn2958, nn2957, 
              nn2956, nn2955} ), 
        .SUM( {\coefcal1_divide_inst1_u126_XORCI_17|SUM_net , dummy_280_, 
              dummy_281_, dummy_282_, dummy_283_, dummy_284_, dummy_285_, dummy_286_, 
              dummy_287_, dummy_288_, dummy_289_, dummy_290_, dummy_291_, dummy_292_, 
              dummy_293_, dummy_294_, dummy_295_, dummy_296_} )
      );
    CS_LUT4_PRIM ii2994 ( .DX(nn2994), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1974_), .F3(dummy_abc_1975_) );
      defparam ii2994.CONFIG_DATA = 16'h9999;
      defparam ii2994.PLACE_LOCATION = "NONE";
      defparam ii2994.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2995 ( .DX(nn2995), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_279_) );
      defparam ii2995.CONFIG_DATA = 16'hA569;
      defparam ii2995.PLACE_LOCATION = "NONE";
      defparam ii2995.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2996 ( .DX(nn2996), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_260_), .F3(dummy_abc_1976_) );
      defparam ii2996.CONFIG_DATA = 16'hA6A6;
      defparam ii2996.PLACE_LOCATION = "NONE";
      defparam ii2996.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2997 ( .DX(nn2997), .F0(dummy_260_), .F1(nn2916), .F2(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ), .F3(dummy_abc_1977_) );
      defparam ii2997.CONFIG_DATA = 16'hD8D8;
      defparam ii2997.PLACE_LOCATION = "NONE";
      defparam ii2997.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2998 ( .DX(nn2998), .F0(nn2917), .F1(dummy_260_), .F2(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ), .F3(dummy_abc_1978_) );
      defparam ii2998.CONFIG_DATA = 16'hB8B8;
      defparam ii2998.PLACE_LOCATION = "NONE";
      defparam ii2998.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2999 ( .DX(nn2999), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1979_), .F3(dummy_abc_1980_) );
      defparam ii2999.CONFIG_DATA = 16'h9999;
      defparam ii2999.PLACE_LOCATION = "NONE";
      defparam ii2999.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3000 ( .DX(nn3000), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_260_) );
      defparam ii3000.CONFIG_DATA = 16'hA569;
      defparam ii3000.PLACE_LOCATION = "NONE";
      defparam ii3000.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3001 ( .DX(nn3001), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_260_), .F2(nn2916), .F3(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ) );
      defparam ii3001.CONFIG_DATA = 16'hA695;
      defparam ii3001.PLACE_LOCATION = "NONE";
      defparam ii3001.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3002 ( .DX(nn3002), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2917), .F2(dummy_260_), .F3(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ) );
      defparam ii3002.CONFIG_DATA = 16'h9A95;
      defparam ii3002.PLACE_LOCATION = "NONE";
      defparam ii3002.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3003 ( .DX(nn3003), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_260_), .F2(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ), .F3(nn2959) );
      defparam ii3003.CONFIG_DATA = 16'hED21;
      defparam ii3003.PLACE_LOCATION = "NONE";
      defparam ii3003.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3004 ( .DX(nn3004), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1981_), .F2(dummy_abc_1982_), .F3(dummy_abc_1983_) );
      defparam ii3004.CONFIG_DATA = 16'h5555;
      defparam ii3004.PLACE_LOCATION = "NONE";
      defparam ii3004.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3005 ( .DX(nn3005), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1984_), .F2(dummy_abc_1985_), .F3(dummy_abc_1986_) );
      defparam ii3005.CONFIG_DATA = 16'h5555;
      defparam ii3005.PLACE_LOCATION = "NONE";
      defparam ii3005.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3006 ( .DX(nn3006), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1987_), .F2(dummy_abc_1988_), .F3(dummy_abc_1989_) );
      defparam ii3006.CONFIG_DATA = 16'h5555;
      defparam ii3006.PLACE_LOCATION = "NONE";
      defparam ii3006.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3007 ( .DX(nn3007), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1990_), .F2(dummy_abc_1991_), .F3(dummy_abc_1992_) );
      defparam ii3007.CONFIG_DATA = 16'h5555;
      defparam ii3007.PLACE_LOCATION = "NONE";
      defparam ii3007.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3008 ( .DX(nn3008), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1993_), .F2(dummy_abc_1994_), .F3(dummy_abc_1995_) );
      defparam ii3008.CONFIG_DATA = 16'h5555;
      defparam ii3008.PLACE_LOCATION = "NONE";
      defparam ii3008.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3009 ( .DX(nn3009), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1996_), .F2(dummy_abc_1997_), .F3(dummy_abc_1998_) );
      defparam ii3009.CONFIG_DATA = 16'h5555;
      defparam ii3009.PLACE_LOCATION = "NONE";
      defparam ii3009.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3010 ( .DX(nn3010), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1999_), .F2(dummy_abc_2000_), .F3(dummy_abc_2001_) );
      defparam ii3010.CONFIG_DATA = 16'h5555;
      defparam ii3010.PLACE_LOCATION = "NONE";
      defparam ii3010.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3011 ( .DX(nn3011), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2002_), .F2(dummy_abc_2003_), .F3(dummy_abc_2004_) );
      defparam ii3011.CONFIG_DATA = 16'h5555;
      defparam ii3011.PLACE_LOCATION = "NONE";
      defparam ii3011.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3012 ( .DX(nn3012), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2005_), .F2(dummy_abc_2006_), .F3(dummy_abc_2007_) );
      defparam ii3012.CONFIG_DATA = 16'h5555;
      defparam ii3012.PLACE_LOCATION = "NONE";
      defparam ii3012.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3013 ( .DX(nn3013), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2008_), .F2(dummy_abc_2009_), .F3(dummy_abc_2010_) );
      defparam ii3013.CONFIG_DATA = 16'h5555;
      defparam ii3013.PLACE_LOCATION = "NONE";
      defparam ii3013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3014 ( .DX(nn3014), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2011_), .F2(dummy_abc_2012_), .F3(dummy_abc_2013_) );
      defparam ii3014.CONFIG_DATA = 16'h5555;
      defparam ii3014.PLACE_LOCATION = "NONE";
      defparam ii3014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3015 ( .DX(nn3015), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2014_), .F2(dummy_abc_2015_), .F3(dummy_abc_2016_) );
      defparam ii3015.CONFIG_DATA = 16'h5555;
      defparam ii3015.PLACE_LOCATION = "NONE";
      defparam ii3015.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_12_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn2954, nn2998, nn2997, nn2996, 
              \coefcal1_xDividend__reg[12]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_144_ ), 
        .DX( {nn3015, nn3014, nn3013, nn3012, nn3011, nn3010, nn3009, nn3008, 
              nn3007, nn3006, nn3005, nn3004, nn3003, nn3002, nn3001, nn3000, 
              nn2999} ), 
        .SUM( {dummy_145_, \coefcal1_divide_inst1_u105_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_14|SUM_net , \coefcal1_divide_inst1_u105_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_12|SUM_net , \coefcal1_divide_inst1_u105_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_10|SUM_net , \coefcal1_divide_inst1_u105_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_8|SUM_net , \coefcal1_divide_inst1_u105_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_6|SUM_net , \coefcal1_divide_inst1_u105_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_4|SUM_net , \coefcal1_divide_inst1_u105_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_2|SUM_net , \coefcal1_divide_inst1_u105_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3035 ( .DX(nn3035), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_279_), .F2(nn2996), .F3(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ) );
      defparam ii3035.CONFIG_DATA = 16'hA695;
      defparam ii3035.PLACE_LOCATION = "NONE";
      defparam ii3035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3036 ( .DX(nn3036), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2997), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ) );
      defparam ii3036.CONFIG_DATA = 16'h9A95;
      defparam ii3036.PLACE_LOCATION = "NONE";
      defparam ii3036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3037 ( .DX(nn3037), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn2998), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ) );
      defparam ii3037.CONFIG_DATA = 16'h9A95;
      defparam ii3037.PLACE_LOCATION = "NONE";
      defparam ii3037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3038 ( .DX(nn3038), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn2954), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_4|SUM_net ) );
      defparam ii3038.CONFIG_DATA = 16'h9A95;
      defparam ii3038.PLACE_LOCATION = "NONE";
      defparam ii3038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3039 ( .DX(nn3039), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2017_), .F2(dummy_abc_2018_), .F3(dummy_abc_2019_) );
      defparam ii3039.CONFIG_DATA = 16'h5555;
      defparam ii3039.PLACE_LOCATION = "NONE";
      defparam ii3039.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3040 ( .DX(nn3040), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2020_), .F2(dummy_abc_2021_), .F3(dummy_abc_2022_) );
      defparam ii3040.CONFIG_DATA = 16'h5555;
      defparam ii3040.PLACE_LOCATION = "NONE";
      defparam ii3040.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3041 ( .DX(nn3041), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2023_), .F2(dummy_abc_2024_), .F3(dummy_abc_2025_) );
      defparam ii3041.CONFIG_DATA = 16'h5555;
      defparam ii3041.PLACE_LOCATION = "NONE";
      defparam ii3041.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3042 ( .DX(nn3042), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2026_), .F2(dummy_abc_2027_), .F3(dummy_abc_2028_) );
      defparam ii3042.CONFIG_DATA = 16'h5555;
      defparam ii3042.PLACE_LOCATION = "NONE";
      defparam ii3042.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3043 ( .DX(nn3043), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2029_), .F2(dummy_abc_2030_), .F3(dummy_abc_2031_) );
      defparam ii3043.CONFIG_DATA = 16'h5555;
      defparam ii3043.PLACE_LOCATION = "NONE";
      defparam ii3043.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3044 ( .DX(nn3044), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2032_), .F2(dummy_abc_2033_), .F3(dummy_abc_2034_) );
      defparam ii3044.CONFIG_DATA = 16'h5555;
      defparam ii3044.PLACE_LOCATION = "NONE";
      defparam ii3044.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3045 ( .DX(nn3045), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2035_), .F2(dummy_abc_2036_), .F3(dummy_abc_2037_) );
      defparam ii3045.CONFIG_DATA = 16'h5555;
      defparam ii3045.PLACE_LOCATION = "NONE";
      defparam ii3045.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3046 ( .DX(nn3046), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2038_), .F2(dummy_abc_2039_), .F3(dummy_abc_2040_) );
      defparam ii3046.CONFIG_DATA = 16'h5555;
      defparam ii3046.PLACE_LOCATION = "NONE";
      defparam ii3046.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3047 ( .DX(nn3047), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2041_), .F2(dummy_abc_2042_), .F3(dummy_abc_2043_) );
      defparam ii3047.CONFIG_DATA = 16'h5555;
      defparam ii3047.PLACE_LOCATION = "NONE";
      defparam ii3047.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3048 ( .DX(nn3048), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2044_), .F2(dummy_abc_2045_), .F3(dummy_abc_2046_) );
      defparam ii3048.CONFIG_DATA = 16'h5555;
      defparam ii3048.PLACE_LOCATION = "NONE";
      defparam ii3048.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3049 ( .DX(nn3049), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2047_), .F2(dummy_abc_2048_), .F3(dummy_abc_2049_) );
      defparam ii3049.CONFIG_DATA = 16'h5555;
      defparam ii3049.PLACE_LOCATION = "NONE";
      defparam ii3049.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3050 ( .DX(nn3050), .F0(dummy_abc_2050_), .F1(dummy_abc_2051_), .F2(dummy_abc_2052_), .F3(dummy_abc_2053_) );
      defparam ii3050.CONFIG_DATA = 16'hFFFF;
      defparam ii3050.PLACE_LOCATION = "NONE";
      defparam ii3050.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_28_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_298_ ), 
        .DX( {nn3050, nn3049, nn3048, nn3047, nn3046, nn3045, nn3044, nn3043, 
              nn3042, nn3041, nn3040, nn3039, nn3038, nn3037, nn3036, nn3035, 
              nn2995, nn2994} ), 
        .SUM( {\coefcal1_divide_inst1_u128_XORCI_17|SUM_net , dummy_299_, 
              dummy_300_, dummy_301_, dummy_302_, dummy_303_, dummy_304_, dummy_305_, 
              dummy_306_, dummy_307_, dummy_308_, dummy_309_, dummy_310_, dummy_311_, 
              dummy_312_, dummy_313_, dummy_314_, dummy_315_} )
      );
    CS_LUT4_PRIM ii3071 ( .DX(nn3071), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_279_), .F3(dummy_abc_2054_) );
      defparam ii3071.CONFIG_DATA = 16'hA6A6;
      defparam ii3071.PLACE_LOCATION = "NONE";
      defparam ii3071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3072 ( .DX(nn3072), .F0(dummy_279_), .F1(nn2996), .F2(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ), .F3(dummy_abc_2055_) );
      defparam ii3072.CONFIG_DATA = 16'hD8D8;
      defparam ii3072.PLACE_LOCATION = "NONE";
      defparam ii3072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3073 ( .DX(nn3073), .F0(nn2997), .F1(dummy_279_), .F2(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ), .F3(dummy_abc_2056_) );
      defparam ii3073.CONFIG_DATA = 16'hB8B8;
      defparam ii3073.PLACE_LOCATION = "NONE";
      defparam ii3073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3074 ( .DX(nn3074), .F0(nn2998), .F1(dummy_279_), .F2(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ), .F3(dummy_abc_2057_) );
      defparam ii3074.CONFIG_DATA = 16'hB8B8;
      defparam ii3074.PLACE_LOCATION = "NONE";
      defparam ii3074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3075 ( .DX(nn3075), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2058_), .F3(dummy_abc_2059_) );
      defparam ii3075.CONFIG_DATA = 16'h9999;
      defparam ii3075.PLACE_LOCATION = "NONE";
      defparam ii3075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3076 ( .DX(nn3076), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_279_) );
      defparam ii3076.CONFIG_DATA = 16'hA569;
      defparam ii3076.PLACE_LOCATION = "NONE";
      defparam ii3076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3077 ( .DX(nn3077), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_279_), .F2(nn2996), .F3(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ) );
      defparam ii3077.CONFIG_DATA = 16'hA695;
      defparam ii3077.PLACE_LOCATION = "NONE";
      defparam ii3077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3078 ( .DX(nn3078), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn2997), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ) );
      defparam ii3078.CONFIG_DATA = 16'h9A95;
      defparam ii3078.PLACE_LOCATION = "NONE";
      defparam ii3078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3079 ( .DX(nn3079), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn2998), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ) );
      defparam ii3079.CONFIG_DATA = 16'h9A95;
      defparam ii3079.PLACE_LOCATION = "NONE";
      defparam ii3079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3080 ( .DX(nn3080), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn2954), .F2(dummy_279_), .F3(\coefcal1_divide_inst1_u105_XORCI_4|SUM_net ) );
      defparam ii3080.CONFIG_DATA = 16'h9A95;
      defparam ii3080.PLACE_LOCATION = "NONE";
      defparam ii3080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3081 ( .DX(nn3081), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2060_), .F2(dummy_abc_2061_), .F3(dummy_abc_2062_) );
      defparam ii3081.CONFIG_DATA = 16'h5555;
      defparam ii3081.PLACE_LOCATION = "NONE";
      defparam ii3081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3082 ( .DX(nn3082), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2063_), .F2(dummy_abc_2064_), .F3(dummy_abc_2065_) );
      defparam ii3082.CONFIG_DATA = 16'h5555;
      defparam ii3082.PLACE_LOCATION = "NONE";
      defparam ii3082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3083 ( .DX(nn3083), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2066_), .F2(dummy_abc_2067_), .F3(dummy_abc_2068_) );
      defparam ii3083.CONFIG_DATA = 16'h5555;
      defparam ii3083.PLACE_LOCATION = "NONE";
      defparam ii3083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3084 ( .DX(nn3084), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2069_), .F2(dummy_abc_2070_), .F3(dummy_abc_2071_) );
      defparam ii3084.CONFIG_DATA = 16'h5555;
      defparam ii3084.PLACE_LOCATION = "NONE";
      defparam ii3084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3085 ( .DX(nn3085), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2072_), .F2(dummy_abc_2073_), .F3(dummy_abc_2074_) );
      defparam ii3085.CONFIG_DATA = 16'h5555;
      defparam ii3085.PLACE_LOCATION = "NONE";
      defparam ii3085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3086 ( .DX(nn3086), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2075_), .F2(dummy_abc_2076_), .F3(dummy_abc_2077_) );
      defparam ii3086.CONFIG_DATA = 16'h5555;
      defparam ii3086.PLACE_LOCATION = "NONE";
      defparam ii3086.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3087 ( .DX(nn3087), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2078_), .F2(dummy_abc_2079_), .F3(dummy_abc_2080_) );
      defparam ii3087.CONFIG_DATA = 16'h5555;
      defparam ii3087.PLACE_LOCATION = "NONE";
      defparam ii3087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3088 ( .DX(nn3088), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2081_), .F2(dummy_abc_2082_), .F3(dummy_abc_2083_) );
      defparam ii3088.CONFIG_DATA = 16'h5555;
      defparam ii3088.PLACE_LOCATION = "NONE";
      defparam ii3088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3089 ( .DX(nn3089), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2084_), .F2(dummy_abc_2085_), .F3(dummy_abc_2086_) );
      defparam ii3089.CONFIG_DATA = 16'h5555;
      defparam ii3089.PLACE_LOCATION = "NONE";
      defparam ii3089.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3090 ( .DX(nn3090), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2087_), .F2(dummy_abc_2088_), .F3(dummy_abc_2089_) );
      defparam ii3090.CONFIG_DATA = 16'h5555;
      defparam ii3090.PLACE_LOCATION = "NONE";
      defparam ii3090.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3091 ( .DX(nn3091), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2090_), .F2(dummy_abc_2091_), .F3(dummy_abc_2092_) );
      defparam ii3091.CONFIG_DATA = 16'h5555;
      defparam ii3091.PLACE_LOCATION = "NONE";
      defparam ii3091.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_13_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn3074, nn3073, nn3072, nn3071, 
              \coefcal1_xDividend__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_146_ ), 
        .DX( {nn3091, nn3090, nn3089, nn3088, nn3087, nn3086, nn3085, nn3084, 
              nn3083, nn3082, nn3081, nn3080, nn3079, nn3078, nn3077, nn3076, 
              nn3075} ), 
        .SUM( {dummy_147_, \coefcal1_divide_inst1_u106_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_14|SUM_net , \coefcal1_divide_inst1_u106_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_12|SUM_net , \coefcal1_divide_inst1_u106_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_10|SUM_net , \coefcal1_divide_inst1_u106_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_8|SUM_net , \coefcal1_divide_inst1_u106_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_6|SUM_net , \coefcal1_divide_inst1_u106_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_4|SUM_net , \coefcal1_divide_inst1_u106_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_2|SUM_net , \coefcal1_divide_inst1_u106_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3111 ( .DX(nn3111), .F0(nn2954), .F1(dummy_279_), .F2(dummy_298_), .F3(\coefcal1_divide_inst1_u106_XORCI_5|SUM_net ) );
      defparam ii3111.CONFIG_DATA = 16'h8A80;
      defparam ii3111.PLACE_LOCATION = "NONE";
      defparam ii3111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3112 ( .DX(nn3112), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2093_), .F3(dummy_abc_2094_) );
      defparam ii3112.CONFIG_DATA = 16'h9999;
      defparam ii3112.PLACE_LOCATION = "NONE";
      defparam ii3112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3113 ( .DX(nn3113), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_298_) );
      defparam ii3113.CONFIG_DATA = 16'hA569;
      defparam ii3113.PLACE_LOCATION = "NONE";
      defparam ii3113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3114 ( .DX(nn3114), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_298_), .F2(nn3071), .F3(\coefcal1_divide_inst1_u106_XORCI_1|SUM_net ) );
      defparam ii3114.CONFIG_DATA = 16'hA695;
      defparam ii3114.PLACE_LOCATION = "NONE";
      defparam ii3114.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3115 ( .DX(nn3115), .F0(nn3072), .F1(dummy_298_), .F2(\coefcal1_divide_inst1_u106_XORCI_2|SUM_net ), .F3(dummy_abc_2095_) );
      defparam ii3115.CONFIG_DATA = 16'hB8B8;
      defparam ii3115.PLACE_LOCATION = "NONE";
      defparam ii3115.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3116 ( .DX(nn3116), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3115), .F2(dummy_abc_2096_), .F3(dummy_abc_2097_) );
      defparam ii3116.CONFIG_DATA = 16'h9999;
      defparam ii3116.PLACE_LOCATION = "NONE";
      defparam ii3116.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3117 ( .DX(nn3117), .F0(nn3073), .F1(dummy_298_), .F2(\coefcal1_divide_inst1_u106_XORCI_3|SUM_net ), .F3(dummy_abc_2098_) );
      defparam ii3117.CONFIG_DATA = 16'hB8B8;
      defparam ii3117.PLACE_LOCATION = "NONE";
      defparam ii3117.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3118 ( .DX(nn3118), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3117), .F2(dummy_abc_2099_), .F3(dummy_abc_2100_) );
      defparam ii3118.CONFIG_DATA = 16'h9999;
      defparam ii3118.PLACE_LOCATION = "NONE";
      defparam ii3118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3119 ( .DX(nn3119), .F0(nn3074), .F1(dummy_298_), .F2(\coefcal1_divide_inst1_u106_XORCI_4|SUM_net ), .F3(dummy_abc_2101_) );
      defparam ii3119.CONFIG_DATA = 16'hB8B8;
      defparam ii3119.PLACE_LOCATION = "NONE";
      defparam ii3119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3120 ( .DX(nn3120), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3119), .F2(dummy_abc_2102_), .F3(dummy_abc_2103_) );
      defparam ii3120.CONFIG_DATA = 16'h9999;
      defparam ii3120.PLACE_LOCATION = "NONE";
      defparam ii3120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3121 ( .DX(nn3121), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3111), .F2(dummy_abc_2104_), .F3(dummy_abc_2105_) );
      defparam ii3121.CONFIG_DATA = 16'h9999;
      defparam ii3121.PLACE_LOCATION = "NONE";
      defparam ii3121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3122 ( .DX(nn3122), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2106_), .F2(dummy_abc_2107_), .F3(dummy_abc_2108_) );
      defparam ii3122.CONFIG_DATA = 16'h5555;
      defparam ii3122.PLACE_LOCATION = "NONE";
      defparam ii3122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3123 ( .DX(nn3123), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2109_), .F2(dummy_abc_2110_), .F3(dummy_abc_2111_) );
      defparam ii3123.CONFIG_DATA = 16'h5555;
      defparam ii3123.PLACE_LOCATION = "NONE";
      defparam ii3123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3124 ( .DX(nn3124), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2112_), .F2(dummy_abc_2113_), .F3(dummy_abc_2114_) );
      defparam ii3124.CONFIG_DATA = 16'h5555;
      defparam ii3124.PLACE_LOCATION = "NONE";
      defparam ii3124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3125 ( .DX(nn3125), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2115_), .F2(dummy_abc_2116_), .F3(dummy_abc_2117_) );
      defparam ii3125.CONFIG_DATA = 16'h5555;
      defparam ii3125.PLACE_LOCATION = "NONE";
      defparam ii3125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3126 ( .DX(nn3126), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2118_), .F2(dummy_abc_2119_), .F3(dummy_abc_2120_) );
      defparam ii3126.CONFIG_DATA = 16'h5555;
      defparam ii3126.PLACE_LOCATION = "NONE";
      defparam ii3126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3127 ( .DX(nn3127), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2121_), .F2(dummy_abc_2122_), .F3(dummy_abc_2123_) );
      defparam ii3127.CONFIG_DATA = 16'h5555;
      defparam ii3127.PLACE_LOCATION = "NONE";
      defparam ii3127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3128 ( .DX(nn3128), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2124_), .F2(dummy_abc_2125_), .F3(dummy_abc_2126_) );
      defparam ii3128.CONFIG_DATA = 16'h5555;
      defparam ii3128.PLACE_LOCATION = "NONE";
      defparam ii3128.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3129 ( .DX(nn3129), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2127_), .F2(dummy_abc_2128_), .F3(dummy_abc_2129_) );
      defparam ii3129.CONFIG_DATA = 16'h5555;
      defparam ii3129.PLACE_LOCATION = "NONE";
      defparam ii3129.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3130 ( .DX(nn3130), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2130_), .F2(dummy_abc_2131_), .F3(dummy_abc_2132_) );
      defparam ii3130.CONFIG_DATA = 16'h5555;
      defparam ii3130.PLACE_LOCATION = "NONE";
      defparam ii3130.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3131 ( .DX(nn3131), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2133_), .F2(dummy_abc_2134_), .F3(dummy_abc_2135_) );
      defparam ii3131.CONFIG_DATA = 16'h5555;
      defparam ii3131.PLACE_LOCATION = "NONE";
      defparam ii3131.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3132 ( .DX(nn3132), .F0(dummy_abc_2136_), .F1(dummy_abc_2137_), .F2(dummy_abc_2138_), .F3(dummy_abc_2139_) );
      defparam ii3132.CONFIG_DATA = 16'hFFFF;
      defparam ii3132.PLACE_LOCATION = "NONE";
      defparam ii3132.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_29_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_317_ ), 
        .DX( {nn3132, nn3131, nn3130, nn3129, nn3128, nn3127, nn3126, nn3125, 
              nn3124, nn3123, nn3122, nn3121, nn3120, nn3118, nn3116, nn3114, 
              nn3113, nn3112} ), 
        .SUM( {\coefcal1_divide_inst1_u130_XORCI_17|SUM_net , dummy_318_, 
              dummy_319_, dummy_320_, dummy_321_, dummy_322_, dummy_323_, dummy_324_, 
              dummy_325_, dummy_326_, dummy_327_, dummy_328_, dummy_329_, dummy_330_, 
              dummy_331_, dummy_332_, dummy_333_, dummy_334_} )
      );
    CS_LUT4_PRIM ii3153 ( .DX(nn3153), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2140_), .F3(dummy_abc_2141_) );
      defparam ii3153.CONFIG_DATA = 16'h9999;
      defparam ii3153.PLACE_LOCATION = "NONE";
      defparam ii3153.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3154 ( .DX(nn3154), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_317_) );
      defparam ii3154.CONFIG_DATA = 16'hA569;
      defparam ii3154.PLACE_LOCATION = "NONE";
      defparam ii3154.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3155 ( .DX(nn3155), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_298_), .F3(dummy_abc_2142_) );
      defparam ii3155.CONFIG_DATA = 16'hA6A6;
      defparam ii3155.PLACE_LOCATION = "NONE";
      defparam ii3155.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3156 ( .DX(nn3156), .F0(dummy_298_), .F1(nn3071), .F2(\coefcal1_divide_inst1_u106_XORCI_1|SUM_net ), .F3(dummy_abc_2143_) );
      defparam ii3156.CONFIG_DATA = 16'hD8D8;
      defparam ii3156.PLACE_LOCATION = "NONE";
      defparam ii3156.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3157 ( .DX(nn3157), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2144_), .F3(dummy_abc_2145_) );
      defparam ii3157.CONFIG_DATA = 16'h9999;
      defparam ii3157.PLACE_LOCATION = "NONE";
      defparam ii3157.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3158 ( .DX(nn3158), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_298_) );
      defparam ii3158.CONFIG_DATA = 16'hA569;
      defparam ii3158.PLACE_LOCATION = "NONE";
      defparam ii3158.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3159 ( .DX(nn3159), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_298_), .F2(nn3071), .F3(\coefcal1_divide_inst1_u106_XORCI_1|SUM_net ) );
      defparam ii3159.CONFIG_DATA = 16'hA695;
      defparam ii3159.PLACE_LOCATION = "NONE";
      defparam ii3159.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3160 ( .DX(nn3160), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3115), .F2(dummy_abc_2146_), .F3(dummy_abc_2147_) );
      defparam ii3160.CONFIG_DATA = 16'h9999;
      defparam ii3160.PLACE_LOCATION = "NONE";
      defparam ii3160.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3161 ( .DX(nn3161), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3117), .F2(dummy_abc_2148_), .F3(dummy_abc_2149_) );
      defparam ii3161.CONFIG_DATA = 16'h9999;
      defparam ii3161.PLACE_LOCATION = "NONE";
      defparam ii3161.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3162 ( .DX(nn3162), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3119), .F2(dummy_abc_2150_), .F3(dummy_abc_2151_) );
      defparam ii3162.CONFIG_DATA = 16'h9999;
      defparam ii3162.PLACE_LOCATION = "NONE";
      defparam ii3162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3163 ( .DX(nn3163), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3111), .F2(dummy_abc_2152_), .F3(dummy_abc_2153_) );
      defparam ii3163.CONFIG_DATA = 16'h9999;
      defparam ii3163.PLACE_LOCATION = "NONE";
      defparam ii3163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3164 ( .DX(nn3164), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2154_), .F2(dummy_abc_2155_), .F3(dummy_abc_2156_) );
      defparam ii3164.CONFIG_DATA = 16'h5555;
      defparam ii3164.PLACE_LOCATION = "NONE";
      defparam ii3164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3165 ( .DX(nn3165), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2157_), .F2(dummy_abc_2158_), .F3(dummy_abc_2159_) );
      defparam ii3165.CONFIG_DATA = 16'h5555;
      defparam ii3165.PLACE_LOCATION = "NONE";
      defparam ii3165.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3166 ( .DX(nn3166), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2160_), .F2(dummy_abc_2161_), .F3(dummy_abc_2162_) );
      defparam ii3166.CONFIG_DATA = 16'h5555;
      defparam ii3166.PLACE_LOCATION = "NONE";
      defparam ii3166.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3167 ( .DX(nn3167), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2163_), .F2(dummy_abc_2164_), .F3(dummy_abc_2165_) );
      defparam ii3167.CONFIG_DATA = 16'h5555;
      defparam ii3167.PLACE_LOCATION = "NONE";
      defparam ii3167.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3168 ( .DX(nn3168), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2166_), .F2(dummy_abc_2167_), .F3(dummy_abc_2168_) );
      defparam ii3168.CONFIG_DATA = 16'h5555;
      defparam ii3168.PLACE_LOCATION = "NONE";
      defparam ii3168.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3169 ( .DX(nn3169), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2169_), .F2(dummy_abc_2170_), .F3(dummy_abc_2171_) );
      defparam ii3169.CONFIG_DATA = 16'h5555;
      defparam ii3169.PLACE_LOCATION = "NONE";
      defparam ii3169.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3170 ( .DX(nn3170), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2172_), .F2(dummy_abc_2173_), .F3(dummy_abc_2174_) );
      defparam ii3170.CONFIG_DATA = 16'h5555;
      defparam ii3170.PLACE_LOCATION = "NONE";
      defparam ii3170.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3171 ( .DX(nn3171), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2175_), .F2(dummy_abc_2176_), .F3(dummy_abc_2177_) );
      defparam ii3171.CONFIG_DATA = 16'h5555;
      defparam ii3171.PLACE_LOCATION = "NONE";
      defparam ii3171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3172 ( .DX(nn3172), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2178_), .F2(dummy_abc_2179_), .F3(dummy_abc_2180_) );
      defparam ii3172.CONFIG_DATA = 16'h5555;
      defparam ii3172.PLACE_LOCATION = "NONE";
      defparam ii3172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3173 ( .DX(nn3173), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2181_), .F2(dummy_abc_2182_), .F3(dummy_abc_2183_) );
      defparam ii3173.CONFIG_DATA = 16'h5555;
      defparam ii3173.PLACE_LOCATION = "NONE";
      defparam ii3173.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_14_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3111, nn3119, nn3117, nn3115, 
              nn3156, nn3155, \coefcal1_xDividend__reg[10]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_148_ ), 
        .DX( {nn3173, nn3172, nn3171, nn3170, nn3169, nn3168, nn3167, nn3166, 
              nn3165, nn3164, nn3163, nn3162, nn3161, nn3160, nn3159, nn3158, 
              nn3157} ), 
        .SUM( {dummy_149_, \coefcal1_divide_inst1_u107_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_14|SUM_net , \coefcal1_divide_inst1_u107_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_12|SUM_net , \coefcal1_divide_inst1_u107_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_10|SUM_net , \coefcal1_divide_inst1_u107_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_8|SUM_net , \coefcal1_divide_inst1_u107_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_6|SUM_net , \coefcal1_divide_inst1_u107_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_4|SUM_net , \coefcal1_divide_inst1_u107_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_2|SUM_net , \coefcal1_divide_inst1_u107_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3193 ( .DX(nn3193), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_317_), .F2(nn3155), .F3(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ) );
      defparam ii3193.CONFIG_DATA = 16'hA695;
      defparam ii3193.PLACE_LOCATION = "NONE";
      defparam ii3193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3194 ( .DX(nn3194), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3156), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ) );
      defparam ii3194.CONFIG_DATA = 16'h9A95;
      defparam ii3194.PLACE_LOCATION = "NONE";
      defparam ii3194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3195 ( .DX(nn3195), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3115), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ) );
      defparam ii3195.CONFIG_DATA = 16'h9A95;
      defparam ii3195.PLACE_LOCATION = "NONE";
      defparam ii3195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3196 ( .DX(nn3196), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3117), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ) );
      defparam ii3196.CONFIG_DATA = 16'h9A95;
      defparam ii3196.PLACE_LOCATION = "NONE";
      defparam ii3196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3197 ( .DX(nn3197), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3119), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ) );
      defparam ii3197.CONFIG_DATA = 16'h9A95;
      defparam ii3197.PLACE_LOCATION = "NONE";
      defparam ii3197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3198 ( .DX(nn3198), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3111), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_6|SUM_net ) );
      defparam ii3198.CONFIG_DATA = 16'h9A95;
      defparam ii3198.PLACE_LOCATION = "NONE";
      defparam ii3198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3199 ( .DX(nn3199), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2184_), .F2(dummy_abc_2185_), .F3(dummy_abc_2186_) );
      defparam ii3199.CONFIG_DATA = 16'h5555;
      defparam ii3199.PLACE_LOCATION = "NONE";
      defparam ii3199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3200 ( .DX(nn3200), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2187_), .F2(dummy_abc_2188_), .F3(dummy_abc_2189_) );
      defparam ii3200.CONFIG_DATA = 16'h5555;
      defparam ii3200.PLACE_LOCATION = "NONE";
      defparam ii3200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3201 ( .DX(nn3201), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2190_), .F2(dummy_abc_2191_), .F3(dummy_abc_2192_) );
      defparam ii3201.CONFIG_DATA = 16'h5555;
      defparam ii3201.PLACE_LOCATION = "NONE";
      defparam ii3201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3202 ( .DX(nn3202), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2193_), .F2(dummy_abc_2194_), .F3(dummy_abc_2195_) );
      defparam ii3202.CONFIG_DATA = 16'h5555;
      defparam ii3202.PLACE_LOCATION = "NONE";
      defparam ii3202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3203 ( .DX(nn3203), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2196_), .F2(dummy_abc_2197_), .F3(dummy_abc_2198_) );
      defparam ii3203.CONFIG_DATA = 16'h5555;
      defparam ii3203.PLACE_LOCATION = "NONE";
      defparam ii3203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3204 ( .DX(nn3204), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2199_), .F2(dummy_abc_2200_), .F3(dummy_abc_2201_) );
      defparam ii3204.CONFIG_DATA = 16'h5555;
      defparam ii3204.PLACE_LOCATION = "NONE";
      defparam ii3204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3205 ( .DX(nn3205), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2202_), .F2(dummy_abc_2203_), .F3(dummy_abc_2204_) );
      defparam ii3205.CONFIG_DATA = 16'h5555;
      defparam ii3205.PLACE_LOCATION = "NONE";
      defparam ii3205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3206 ( .DX(nn3206), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2205_), .F2(dummy_abc_2206_), .F3(dummy_abc_2207_) );
      defparam ii3206.CONFIG_DATA = 16'h5555;
      defparam ii3206.PLACE_LOCATION = "NONE";
      defparam ii3206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3207 ( .DX(nn3207), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2208_), .F2(dummy_abc_2209_), .F3(dummy_abc_2210_) );
      defparam ii3207.CONFIG_DATA = 16'h5555;
      defparam ii3207.PLACE_LOCATION = "NONE";
      defparam ii3207.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3208 ( .DX(nn3208), .F0(dummy_abc_2211_), .F1(dummy_abc_2212_), .F2(dummy_abc_2213_), .F3(dummy_abc_2214_) );
      defparam ii3208.CONFIG_DATA = 16'hFFFF;
      defparam ii3208.PLACE_LOCATION = "NONE";
      defparam ii3208.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_30_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_336_ ), 
        .DX( {nn3208, nn3207, nn3206, nn3205, nn3204, nn3203, nn3202, nn3201, 
              nn3200, nn3199, nn3198, nn3197, nn3196, nn3195, nn3194, nn3193, 
              nn3154, nn3153} ), 
        .SUM( {\coefcal1_divide_inst1_u132_XORCI_17|SUM_net , dummy_337_, 
              dummy_338_, dummy_339_, dummy_340_, dummy_341_, dummy_342_, dummy_343_, 
              dummy_344_, dummy_345_, dummy_346_, dummy_347_, dummy_348_, dummy_349_, 
              dummy_350_, dummy_351_, dummy_352_, dummy_353_} )
      );
    CS_LUT4_PRIM ii3229 ( .DX(nn3229), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_317_), .F3(dummy_abc_2215_) );
      defparam ii3229.CONFIG_DATA = 16'hA6A6;
      defparam ii3229.PLACE_LOCATION = "NONE";
      defparam ii3229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3230 ( .DX(nn3230), .F0(dummy_317_), .F1(nn3155), .F2(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ), .F3(dummy_abc_2216_) );
      defparam ii3230.CONFIG_DATA = 16'hD8D8;
      defparam ii3230.PLACE_LOCATION = "NONE";
      defparam ii3230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3231 ( .DX(nn3231), .F0(nn3156), .F1(dummy_317_), .F2(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ), .F3(dummy_abc_2217_) );
      defparam ii3231.CONFIG_DATA = 16'hB8B8;
      defparam ii3231.PLACE_LOCATION = "NONE";
      defparam ii3231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3232 ( .DX(nn3232), .F0(nn3115), .F1(dummy_317_), .F2(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ), .F3(dummy_abc_2218_) );
      defparam ii3232.CONFIG_DATA = 16'hB8B8;
      defparam ii3232.PLACE_LOCATION = "NONE";
      defparam ii3232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3233 ( .DX(nn3233), .F0(nn3117), .F1(dummy_317_), .F2(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ), .F3(dummy_abc_2219_) );
      defparam ii3233.CONFIG_DATA = 16'hB8B8;
      defparam ii3233.PLACE_LOCATION = "NONE";
      defparam ii3233.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3234 ( .DX(nn3234), .F0(nn3119), .F1(dummy_317_), .F2(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ), .F3(dummy_abc_2220_) );
      defparam ii3234.CONFIG_DATA = 16'hB8B8;
      defparam ii3234.PLACE_LOCATION = "NONE";
      defparam ii3234.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3235 ( .DX(nn3235), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2221_), .F3(dummy_abc_2222_) );
      defparam ii3235.CONFIG_DATA = 16'h9999;
      defparam ii3235.PLACE_LOCATION = "NONE";
      defparam ii3235.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3236 ( .DX(nn3236), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_317_) );
      defparam ii3236.CONFIG_DATA = 16'hA569;
      defparam ii3236.PLACE_LOCATION = "NONE";
      defparam ii3236.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3237 ( .DX(nn3237), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_317_), .F2(nn3155), .F3(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ) );
      defparam ii3237.CONFIG_DATA = 16'hA695;
      defparam ii3237.PLACE_LOCATION = "NONE";
      defparam ii3237.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3238 ( .DX(nn3238), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3156), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ) );
      defparam ii3238.CONFIG_DATA = 16'h9A95;
      defparam ii3238.PLACE_LOCATION = "NONE";
      defparam ii3238.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3239 ( .DX(nn3239), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3115), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ) );
      defparam ii3239.CONFIG_DATA = 16'h9A95;
      defparam ii3239.PLACE_LOCATION = "NONE";
      defparam ii3239.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3240 ( .DX(nn3240), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3117), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ) );
      defparam ii3240.CONFIG_DATA = 16'h9A95;
      defparam ii3240.PLACE_LOCATION = "NONE";
      defparam ii3240.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3241 ( .DX(nn3241), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3119), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ) );
      defparam ii3241.CONFIG_DATA = 16'h9A95;
      defparam ii3241.PLACE_LOCATION = "NONE";
      defparam ii3241.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3242 ( .DX(nn3242), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3111), .F2(dummy_317_), .F3(\coefcal1_divide_inst1_u107_XORCI_6|SUM_net ) );
      defparam ii3242.CONFIG_DATA = 16'h9A95;
      defparam ii3242.PLACE_LOCATION = "NONE";
      defparam ii3242.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3243 ( .DX(nn3243), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2223_), .F2(dummy_abc_2224_), .F3(dummy_abc_2225_) );
      defparam ii3243.CONFIG_DATA = 16'h5555;
      defparam ii3243.PLACE_LOCATION = "NONE";
      defparam ii3243.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3244 ( .DX(nn3244), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2226_), .F2(dummy_abc_2227_), .F3(dummy_abc_2228_) );
      defparam ii3244.CONFIG_DATA = 16'h5555;
      defparam ii3244.PLACE_LOCATION = "NONE";
      defparam ii3244.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3245 ( .DX(nn3245), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2229_), .F2(dummy_abc_2230_), .F3(dummy_abc_2231_) );
      defparam ii3245.CONFIG_DATA = 16'h5555;
      defparam ii3245.PLACE_LOCATION = "NONE";
      defparam ii3245.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3246 ( .DX(nn3246), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2232_), .F2(dummy_abc_2233_), .F3(dummy_abc_2234_) );
      defparam ii3246.CONFIG_DATA = 16'h5555;
      defparam ii3246.PLACE_LOCATION = "NONE";
      defparam ii3246.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3247 ( .DX(nn3247), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2235_), .F2(dummy_abc_2236_), .F3(dummy_abc_2237_) );
      defparam ii3247.CONFIG_DATA = 16'h5555;
      defparam ii3247.PLACE_LOCATION = "NONE";
      defparam ii3247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3248 ( .DX(nn3248), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2238_), .F2(dummy_abc_2239_), .F3(dummy_abc_2240_) );
      defparam ii3248.CONFIG_DATA = 16'h5555;
      defparam ii3248.PLACE_LOCATION = "NONE";
      defparam ii3248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3249 ( .DX(nn3249), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2241_), .F2(dummy_abc_2242_), .F3(dummy_abc_2243_) );
      defparam ii3249.CONFIG_DATA = 16'h5555;
      defparam ii3249.PLACE_LOCATION = "NONE";
      defparam ii3249.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3250 ( .DX(nn3250), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2244_), .F2(dummy_abc_2245_), .F3(dummy_abc_2246_) );
      defparam ii3250.CONFIG_DATA = 16'h5555;
      defparam ii3250.PLACE_LOCATION = "NONE";
      defparam ii3250.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3251 ( .DX(nn3251), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2247_), .F2(dummy_abc_2248_), .F3(dummy_abc_2249_) );
      defparam ii3251.CONFIG_DATA = 16'h5555;
      defparam ii3251.PLACE_LOCATION = "NONE";
      defparam ii3251.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_15_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3234, nn3233, nn3232, nn3231, 
              nn3230, nn3229, \coefcal1_xDividend__reg[9]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_150_ ), 
        .DX( {nn3251, nn3250, nn3249, nn3248, nn3247, nn3246, nn3245, nn3244, 
              nn3243, nn3242, nn3241, nn3240, nn3239, nn3238, nn3237, nn3236, 
              nn3235} ), 
        .SUM( {dummy_151_, \coefcal1_divide_inst1_u108_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_14|SUM_net , \coefcal1_divide_inst1_u108_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_12|SUM_net , \coefcal1_divide_inst1_u108_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_10|SUM_net , \coefcal1_divide_inst1_u108_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_8|SUM_net , \coefcal1_divide_inst1_u108_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_6|SUM_net , \coefcal1_divide_inst1_u108_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_4|SUM_net , \coefcal1_divide_inst1_u108_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_2|SUM_net , \coefcal1_divide_inst1_u108_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3271 ( .DX(nn3271), .F0(nn3111), .F1(dummy_317_), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ) );
      defparam ii3271.CONFIG_DATA = 16'h8F80;
      defparam ii3271.PLACE_LOCATION = "NONE";
      defparam ii3271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3272 ( .DX(nn3272), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2250_), .F3(dummy_abc_2251_) );
      defparam ii3272.CONFIG_DATA = 16'h9999;
      defparam ii3272.PLACE_LOCATION = "NONE";
      defparam ii3272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3273 ( .DX(nn3273), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_336_) );
      defparam ii3273.CONFIG_DATA = 16'hA569;
      defparam ii3273.PLACE_LOCATION = "NONE";
      defparam ii3273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3274 ( .DX(nn3274), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_336_), .F2(nn3229), .F3(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ) );
      defparam ii3274.CONFIG_DATA = 16'hA695;
      defparam ii3274.PLACE_LOCATION = "NONE";
      defparam ii3274.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3275 ( .DX(nn3275), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3230), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ) );
      defparam ii3275.CONFIG_DATA = 16'h9A95;
      defparam ii3275.PLACE_LOCATION = "NONE";
      defparam ii3275.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3276 ( .DX(nn3276), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3231), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ) );
      defparam ii3276.CONFIG_DATA = 16'h9A95;
      defparam ii3276.PLACE_LOCATION = "NONE";
      defparam ii3276.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3277 ( .DX(nn3277), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3232), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ) );
      defparam ii3277.CONFIG_DATA = 16'h9A95;
      defparam ii3277.PLACE_LOCATION = "NONE";
      defparam ii3277.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3278 ( .DX(nn3278), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3233), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ) );
      defparam ii3278.CONFIG_DATA = 16'h9A95;
      defparam ii3278.PLACE_LOCATION = "NONE";
      defparam ii3278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3279 ( .DX(nn3279), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3234), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ) );
      defparam ii3279.CONFIG_DATA = 16'h9A95;
      defparam ii3279.PLACE_LOCATION = "NONE";
      defparam ii3279.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3280 ( .DX(nn3280), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3111), .F2(dummy_317_), .F3(dummy_abc_2252_) );
      defparam ii3280.CONFIG_DATA = 16'h9595;
      defparam ii3280.PLACE_LOCATION = "NONE";
      defparam ii3280.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3281 ( .DX(nn3281), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ), .F3(nn3280) );
      defparam ii3281.CONFIG_DATA = 16'hCD01;
      defparam ii3281.PLACE_LOCATION = "NONE";
      defparam ii3281.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3282 ( .DX(nn3282), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2253_), .F2(dummy_abc_2254_), .F3(dummy_abc_2255_) );
      defparam ii3282.CONFIG_DATA = 16'h5555;
      defparam ii3282.PLACE_LOCATION = "NONE";
      defparam ii3282.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3283 ( .DX(nn3283), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2256_), .F2(dummy_abc_2257_), .F3(dummy_abc_2258_) );
      defparam ii3283.CONFIG_DATA = 16'h5555;
      defparam ii3283.PLACE_LOCATION = "NONE";
      defparam ii3283.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3284 ( .DX(nn3284), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2259_), .F2(dummy_abc_2260_), .F3(dummy_abc_2261_) );
      defparam ii3284.CONFIG_DATA = 16'h5555;
      defparam ii3284.PLACE_LOCATION = "NONE";
      defparam ii3284.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3285 ( .DX(nn3285), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2262_), .F2(dummy_abc_2263_), .F3(dummy_abc_2264_) );
      defparam ii3285.CONFIG_DATA = 16'h5555;
      defparam ii3285.PLACE_LOCATION = "NONE";
      defparam ii3285.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3286 ( .DX(nn3286), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2265_), .F2(dummy_abc_2266_), .F3(dummy_abc_2267_) );
      defparam ii3286.CONFIG_DATA = 16'h5555;
      defparam ii3286.PLACE_LOCATION = "NONE";
      defparam ii3286.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3287 ( .DX(nn3287), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2268_), .F2(dummy_abc_2269_), .F3(dummy_abc_2270_) );
      defparam ii3287.CONFIG_DATA = 16'h5555;
      defparam ii3287.PLACE_LOCATION = "NONE";
      defparam ii3287.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3288 ( .DX(nn3288), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2271_), .F2(dummy_abc_2272_), .F3(dummy_abc_2273_) );
      defparam ii3288.CONFIG_DATA = 16'h5555;
      defparam ii3288.PLACE_LOCATION = "NONE";
      defparam ii3288.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3289 ( .DX(nn3289), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2274_), .F2(dummy_abc_2275_), .F3(dummy_abc_2276_) );
      defparam ii3289.CONFIG_DATA = 16'h5555;
      defparam ii3289.PLACE_LOCATION = "NONE";
      defparam ii3289.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3290 ( .DX(nn3290), .F0(dummy_abc_2277_), .F1(dummy_abc_2278_), .F2(dummy_abc_2279_), .F3(dummy_abc_2280_) );
      defparam ii3290.CONFIG_DATA = 16'hFFFF;
      defparam ii3290.PLACE_LOCATION = "NONE";
      defparam ii3290.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_31_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_355_ ), 
        .DX( {nn3290, nn3289, nn3288, nn3287, nn3286, nn3285, nn3284, nn3283, 
              nn3282, nn3281, nn3279, nn3278, nn3277, nn3276, nn3275, nn3274, 
              nn3273, nn3272} ), 
        .SUM( {\coefcal1_divide_inst1_u134_XORCI_17|SUM_net , dummy_356_, 
              dummy_357_, dummy_358_, dummy_359_, dummy_360_, dummy_361_, dummy_362_, 
              dummy_363_, dummy_364_, dummy_365_, dummy_366_, dummy_367_, dummy_368_, 
              dummy_369_, dummy_370_, dummy_371_, dummy_372_} )
      );
    CS_LUT4_PRIM ii3311 ( .DX(nn3311), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_336_), .F3(dummy_abc_2281_) );
      defparam ii3311.CONFIG_DATA = 16'hA6A6;
      defparam ii3311.PLACE_LOCATION = "NONE";
      defparam ii3311.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3312 ( .DX(nn3312), .F0(dummy_336_), .F1(nn3229), .F2(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ), .F3(dummy_abc_2282_) );
      defparam ii3312.CONFIG_DATA = 16'hD8D8;
      defparam ii3312.PLACE_LOCATION = "NONE";
      defparam ii3312.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3313 ( .DX(nn3313), .F0(nn3230), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ), .F3(dummy_abc_2283_) );
      defparam ii3313.CONFIG_DATA = 16'hB8B8;
      defparam ii3313.PLACE_LOCATION = "NONE";
      defparam ii3313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3314 ( .DX(nn3314), .F0(nn3231), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ), .F3(dummy_abc_2284_) );
      defparam ii3314.CONFIG_DATA = 16'hB8B8;
      defparam ii3314.PLACE_LOCATION = "NONE";
      defparam ii3314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3315 ( .DX(nn3315), .F0(nn3232), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ), .F3(dummy_abc_2285_) );
      defparam ii3315.CONFIG_DATA = 16'hB8B8;
      defparam ii3315.PLACE_LOCATION = "NONE";
      defparam ii3315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3316 ( .DX(nn3316), .F0(nn3233), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ), .F3(dummy_abc_2286_) );
      defparam ii3316.CONFIG_DATA = 16'hB8B8;
      defparam ii3316.PLACE_LOCATION = "NONE";
      defparam ii3316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3317 ( .DX(nn3317), .F0(nn3234), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ), .F3(dummy_abc_2287_) );
      defparam ii3317.CONFIG_DATA = 16'hB8B8;
      defparam ii3317.PLACE_LOCATION = "NONE";
      defparam ii3317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3318 ( .DX(nn3318), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2288_), .F3(dummy_abc_2289_) );
      defparam ii3318.CONFIG_DATA = 16'h9999;
      defparam ii3318.PLACE_LOCATION = "NONE";
      defparam ii3318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3319 ( .DX(nn3319), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_336_) );
      defparam ii3319.CONFIG_DATA = 16'hA569;
      defparam ii3319.PLACE_LOCATION = "NONE";
      defparam ii3319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3320 ( .DX(nn3320), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_336_), .F2(nn3229), .F3(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ) );
      defparam ii3320.CONFIG_DATA = 16'hA695;
      defparam ii3320.PLACE_LOCATION = "NONE";
      defparam ii3320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3321 ( .DX(nn3321), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3230), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ) );
      defparam ii3321.CONFIG_DATA = 16'h9A95;
      defparam ii3321.PLACE_LOCATION = "NONE";
      defparam ii3321.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3322 ( .DX(nn3322), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3231), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ) );
      defparam ii3322.CONFIG_DATA = 16'h9A95;
      defparam ii3322.PLACE_LOCATION = "NONE";
      defparam ii3322.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3323 ( .DX(nn3323), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3232), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ) );
      defparam ii3323.CONFIG_DATA = 16'h9A95;
      defparam ii3323.PLACE_LOCATION = "NONE";
      defparam ii3323.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3324 ( .DX(nn3324), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3233), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ) );
      defparam ii3324.CONFIG_DATA = 16'h9A95;
      defparam ii3324.PLACE_LOCATION = "NONE";
      defparam ii3324.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3325 ( .DX(nn3325), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3234), .F2(dummy_336_), .F3(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ) );
      defparam ii3325.CONFIG_DATA = 16'h9A95;
      defparam ii3325.PLACE_LOCATION = "NONE";
      defparam ii3325.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3326 ( .DX(nn3326), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_336_), .F2(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ), .F3(nn3280) );
      defparam ii3326.CONFIG_DATA = 16'hCD01;
      defparam ii3326.PLACE_LOCATION = "NONE";
      defparam ii3326.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3327 ( .DX(nn3327), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2290_), .F2(dummy_abc_2291_), .F3(dummy_abc_2292_) );
      defparam ii3327.CONFIG_DATA = 16'h5555;
      defparam ii3327.PLACE_LOCATION = "NONE";
      defparam ii3327.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3328 ( .DX(nn3328), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2293_), .F2(dummy_abc_2294_), .F3(dummy_abc_2295_) );
      defparam ii3328.CONFIG_DATA = 16'h5555;
      defparam ii3328.PLACE_LOCATION = "NONE";
      defparam ii3328.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3329 ( .DX(nn3329), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2296_), .F2(dummy_abc_2297_), .F3(dummy_abc_2298_) );
      defparam ii3329.CONFIG_DATA = 16'h5555;
      defparam ii3329.PLACE_LOCATION = "NONE";
      defparam ii3329.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3330 ( .DX(nn3330), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2299_), .F2(dummy_abc_2300_), .F3(dummy_abc_2301_) );
      defparam ii3330.CONFIG_DATA = 16'h5555;
      defparam ii3330.PLACE_LOCATION = "NONE";
      defparam ii3330.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3331 ( .DX(nn3331), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2302_), .F2(dummy_abc_2303_), .F3(dummy_abc_2304_) );
      defparam ii3331.CONFIG_DATA = 16'h5555;
      defparam ii3331.PLACE_LOCATION = "NONE";
      defparam ii3331.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3332 ( .DX(nn3332), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2305_), .F2(dummy_abc_2306_), .F3(dummy_abc_2307_) );
      defparam ii3332.CONFIG_DATA = 16'h5555;
      defparam ii3332.PLACE_LOCATION = "NONE";
      defparam ii3332.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3333 ( .DX(nn3333), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2308_), .F2(dummy_abc_2309_), .F3(dummy_abc_2310_) );
      defparam ii3333.CONFIG_DATA = 16'h5555;
      defparam ii3333.PLACE_LOCATION = "NONE";
      defparam ii3333.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3334 ( .DX(nn3334), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2311_), .F2(dummy_abc_2312_), .F3(dummy_abc_2313_) );
      defparam ii3334.CONFIG_DATA = 16'h5555;
      defparam ii3334.PLACE_LOCATION = "NONE";
      defparam ii3334.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_16_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3271, 
              nn3317, nn3316, nn3315, nn3314, nn3313, nn3312, nn3311, 
              \coefcal1_xDividend__reg[8]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_152_ ), 
        .DX( {nn3334, nn3333, nn3332, nn3331, nn3330, nn3329, nn3328, nn3327, 
              nn3326, nn3325, nn3324, nn3323, nn3322, nn3321, nn3320, nn3319, 
              nn3318} ), 
        .SUM( {dummy_153_, \coefcal1_divide_inst1_u109_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_14|SUM_net , \coefcal1_divide_inst1_u109_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_12|SUM_net , \coefcal1_divide_inst1_u109_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_10|SUM_net , \coefcal1_divide_inst1_u109_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_8|SUM_net , \coefcal1_divide_inst1_u109_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_6|SUM_net , \coefcal1_divide_inst1_u109_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_4|SUM_net , \coefcal1_divide_inst1_u109_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_2|SUM_net , \coefcal1_divide_inst1_u109_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3354 ( .DX(nn3354), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2314_), .F3(dummy_abc_2315_) );
      defparam ii3354.CONFIG_DATA = 16'h9999;
      defparam ii3354.PLACE_LOCATION = "NONE";
      defparam ii3354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3355 ( .DX(nn3355), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_355_) );
      defparam ii3355.CONFIG_DATA = 16'hA569;
      defparam ii3355.PLACE_LOCATION = "NONE";
      defparam ii3355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3356 ( .DX(nn3356), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_355_), .F2(nn3311), .F3(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ) );
      defparam ii3356.CONFIG_DATA = 16'hA695;
      defparam ii3356.PLACE_LOCATION = "NONE";
      defparam ii3356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3357 ( .DX(nn3357), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3312), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ) );
      defparam ii3357.CONFIG_DATA = 16'h9A95;
      defparam ii3357.PLACE_LOCATION = "NONE";
      defparam ii3357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3358 ( .DX(nn3358), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3313), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ) );
      defparam ii3358.CONFIG_DATA = 16'h9A95;
      defparam ii3358.PLACE_LOCATION = "NONE";
      defparam ii3358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3359 ( .DX(nn3359), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3314), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ) );
      defparam ii3359.CONFIG_DATA = 16'h9A95;
      defparam ii3359.PLACE_LOCATION = "NONE";
      defparam ii3359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3360 ( .DX(nn3360), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3315), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ) );
      defparam ii3360.CONFIG_DATA = 16'h9A95;
      defparam ii3360.PLACE_LOCATION = "NONE";
      defparam ii3360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3361 ( .DX(nn3361), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3316), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ) );
      defparam ii3361.CONFIG_DATA = 16'h9A95;
      defparam ii3361.PLACE_LOCATION = "NONE";
      defparam ii3361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3362 ( .DX(nn3362), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3317), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ) );
      defparam ii3362.CONFIG_DATA = 16'h9A95;
      defparam ii3362.PLACE_LOCATION = "NONE";
      defparam ii3362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3363 ( .DX(nn3363), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3271), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ) );
      defparam ii3363.CONFIG_DATA = 16'h9995;
      defparam ii3363.PLACE_LOCATION = "NONE";
      defparam ii3363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3364 ( .DX(nn3364), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2316_), .F2(dummy_abc_2317_), .F3(dummy_abc_2318_) );
      defparam ii3364.CONFIG_DATA = 16'h5555;
      defparam ii3364.PLACE_LOCATION = "NONE";
      defparam ii3364.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3365 ( .DX(nn3365), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2319_), .F2(dummy_abc_2320_), .F3(dummy_abc_2321_) );
      defparam ii3365.CONFIG_DATA = 16'h5555;
      defparam ii3365.PLACE_LOCATION = "NONE";
      defparam ii3365.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3366 ( .DX(nn3366), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2322_), .F2(dummy_abc_2323_), .F3(dummy_abc_2324_) );
      defparam ii3366.CONFIG_DATA = 16'h5555;
      defparam ii3366.PLACE_LOCATION = "NONE";
      defparam ii3366.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3367 ( .DX(nn3367), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2325_), .F2(dummy_abc_2326_), .F3(dummy_abc_2327_) );
      defparam ii3367.CONFIG_DATA = 16'h5555;
      defparam ii3367.PLACE_LOCATION = "NONE";
      defparam ii3367.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3368 ( .DX(nn3368), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2328_), .F2(dummy_abc_2329_), .F3(dummy_abc_2330_) );
      defparam ii3368.CONFIG_DATA = 16'h5555;
      defparam ii3368.PLACE_LOCATION = "NONE";
      defparam ii3368.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3369 ( .DX(nn3369), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2331_), .F2(dummy_abc_2332_), .F3(dummy_abc_2333_) );
      defparam ii3369.CONFIG_DATA = 16'h5555;
      defparam ii3369.PLACE_LOCATION = "NONE";
      defparam ii3369.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3370 ( .DX(nn3370), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2334_), .F2(dummy_abc_2335_), .F3(dummy_abc_2336_) );
      defparam ii3370.CONFIG_DATA = 16'h5555;
      defparam ii3370.PLACE_LOCATION = "NONE";
      defparam ii3370.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3371 ( .DX(nn3371), .F0(dummy_abc_2337_), .F1(dummy_abc_2338_), .F2(dummy_abc_2339_), .F3(dummy_abc_2340_) );
      defparam ii3371.CONFIG_DATA = 16'hFFFF;
      defparam ii3371.PLACE_LOCATION = "NONE";
      defparam ii3371.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_32_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_374_ ), 
        .DX( {nn3371, nn3370, nn3369, nn3368, nn3367, nn3366, nn3365, nn3364, 
              nn3363, nn3362, nn3361, nn3360, nn3359, nn3358, nn3357, nn3356, 
              nn3355, nn3354} ), 
        .SUM( {\coefcal1_divide_inst1_u136_XORCI_17|SUM_net , dummy_375_, 
              dummy_376_, dummy_377_, dummy_378_, dummy_379_, dummy_380_, dummy_381_, 
              dummy_382_, dummy_383_, dummy_384_, dummy_385_, dummy_386_, dummy_387_, 
              dummy_388_, dummy_389_, dummy_390_, dummy_391_} )
      );
    CS_LUT4_PRIM ii3392 ( .DX(nn3392), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_355_), .F3(dummy_abc_2341_) );
      defparam ii3392.CONFIG_DATA = 16'hA6A6;
      defparam ii3392.PLACE_LOCATION = "NONE";
      defparam ii3392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3393 ( .DX(nn3393), .F0(dummy_355_), .F1(nn3311), .F2(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ), .F3(dummy_abc_2342_) );
      defparam ii3393.CONFIG_DATA = 16'hD8D8;
      defparam ii3393.PLACE_LOCATION = "NONE";
      defparam ii3393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3394 ( .DX(nn3394), .F0(nn3312), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ), .F3(dummy_abc_2343_) );
      defparam ii3394.CONFIG_DATA = 16'hB8B8;
      defparam ii3394.PLACE_LOCATION = "NONE";
      defparam ii3394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3395 ( .DX(nn3395), .F0(nn3313), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ), .F3(dummy_abc_2344_) );
      defparam ii3395.CONFIG_DATA = 16'hB8B8;
      defparam ii3395.PLACE_LOCATION = "NONE";
      defparam ii3395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3396 ( .DX(nn3396), .F0(nn3314), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ), .F3(dummy_abc_2345_) );
      defparam ii3396.CONFIG_DATA = 16'hB8B8;
      defparam ii3396.PLACE_LOCATION = "NONE";
      defparam ii3396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3397 ( .DX(nn3397), .F0(nn3315), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ), .F3(dummy_abc_2346_) );
      defparam ii3397.CONFIG_DATA = 16'hB8B8;
      defparam ii3397.PLACE_LOCATION = "NONE";
      defparam ii3397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3398 ( .DX(nn3398), .F0(nn3316), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ), .F3(dummy_abc_2347_) );
      defparam ii3398.CONFIG_DATA = 16'hB8B8;
      defparam ii3398.PLACE_LOCATION = "NONE";
      defparam ii3398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3399 ( .DX(nn3399), .F0(nn3317), .F1(dummy_355_), .F2(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ), .F3(dummy_abc_2348_) );
      defparam ii3399.CONFIG_DATA = 16'hB8B8;
      defparam ii3399.PLACE_LOCATION = "NONE";
      defparam ii3399.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3400 ( .DX(nn3400), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2349_), .F3(dummy_abc_2350_) );
      defparam ii3400.CONFIG_DATA = 16'h9999;
      defparam ii3400.PLACE_LOCATION = "NONE";
      defparam ii3400.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3401 ( .DX(nn3401), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_355_) );
      defparam ii3401.CONFIG_DATA = 16'hA569;
      defparam ii3401.PLACE_LOCATION = "NONE";
      defparam ii3401.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3402 ( .DX(nn3402), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_355_), .F2(nn3311), .F3(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ) );
      defparam ii3402.CONFIG_DATA = 16'hA695;
      defparam ii3402.PLACE_LOCATION = "NONE";
      defparam ii3402.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3403 ( .DX(nn3403), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3312), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ) );
      defparam ii3403.CONFIG_DATA = 16'h9A95;
      defparam ii3403.PLACE_LOCATION = "NONE";
      defparam ii3403.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3404 ( .DX(nn3404), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3313), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ) );
      defparam ii3404.CONFIG_DATA = 16'h9A95;
      defparam ii3404.PLACE_LOCATION = "NONE";
      defparam ii3404.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3405 ( .DX(nn3405), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3314), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ) );
      defparam ii3405.CONFIG_DATA = 16'h9A95;
      defparam ii3405.PLACE_LOCATION = "NONE";
      defparam ii3405.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3406 ( .DX(nn3406), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3315), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ) );
      defparam ii3406.CONFIG_DATA = 16'h9A95;
      defparam ii3406.PLACE_LOCATION = "NONE";
      defparam ii3406.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3407 ( .DX(nn3407), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3316), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ) );
      defparam ii3407.CONFIG_DATA = 16'h9A95;
      defparam ii3407.PLACE_LOCATION = "NONE";
      defparam ii3407.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3408 ( .DX(nn3408), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3317), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ) );
      defparam ii3408.CONFIG_DATA = 16'h9A95;
      defparam ii3408.PLACE_LOCATION = "NONE";
      defparam ii3408.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3409 ( .DX(nn3409), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3271), .F2(dummy_355_), .F3(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ) );
      defparam ii3409.CONFIG_DATA = 16'h9995;
      defparam ii3409.PLACE_LOCATION = "NONE";
      defparam ii3409.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3410 ( .DX(nn3410), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2351_), .F2(dummy_abc_2352_), .F3(dummy_abc_2353_) );
      defparam ii3410.CONFIG_DATA = 16'h5555;
      defparam ii3410.PLACE_LOCATION = "NONE";
      defparam ii3410.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3411 ( .DX(nn3411), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2354_), .F2(dummy_abc_2355_), .F3(dummy_abc_2356_) );
      defparam ii3411.CONFIG_DATA = 16'h5555;
      defparam ii3411.PLACE_LOCATION = "NONE";
      defparam ii3411.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3412 ( .DX(nn3412), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2357_), .F2(dummy_abc_2358_), .F3(dummy_abc_2359_) );
      defparam ii3412.CONFIG_DATA = 16'h5555;
      defparam ii3412.PLACE_LOCATION = "NONE";
      defparam ii3412.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3413 ( .DX(nn3413), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2360_), .F2(dummy_abc_2361_), .F3(dummy_abc_2362_) );
      defparam ii3413.CONFIG_DATA = 16'h5555;
      defparam ii3413.PLACE_LOCATION = "NONE";
      defparam ii3413.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3414 ( .DX(nn3414), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2363_), .F2(dummy_abc_2364_), .F3(dummy_abc_2365_) );
      defparam ii3414.CONFIG_DATA = 16'h5555;
      defparam ii3414.PLACE_LOCATION = "NONE";
      defparam ii3414.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3415 ( .DX(nn3415), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2366_), .F2(dummy_abc_2367_), .F3(dummy_abc_2368_) );
      defparam ii3415.CONFIG_DATA = 16'h5555;
      defparam ii3415.PLACE_LOCATION = "NONE";
      defparam ii3415.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3416 ( .DX(nn3416), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2369_), .F2(dummy_abc_2370_), .F3(dummy_abc_2371_) );
      defparam ii3416.CONFIG_DATA = 16'h5555;
      defparam ii3416.PLACE_LOCATION = "NONE";
      defparam ii3416.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_17_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3399, 
              nn3398, nn3397, nn3396, nn3395, nn3394, nn3393, nn3392, 
              \coefcal1_xDividend__reg[7]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_154_ ), 
        .DX( {nn3416, nn3415, nn3414, nn3413, nn3412, nn3411, nn3410, nn3409, 
              nn3408, nn3407, nn3406, nn3405, nn3404, nn3403, nn3402, nn3401, 
              nn3400} ), 
        .SUM( {dummy_155_, \coefcal1_divide_inst1_u110_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_14|SUM_net , \coefcal1_divide_inst1_u110_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_12|SUM_net , \coefcal1_divide_inst1_u110_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_10|SUM_net , \coefcal1_divide_inst1_u110_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_8|SUM_net , \coefcal1_divide_inst1_u110_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_6|SUM_net , \coefcal1_divide_inst1_u110_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_4|SUM_net , \coefcal1_divide_inst1_u110_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_2|SUM_net , \coefcal1_divide_inst1_u110_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3436 ( .DX(nn3436), .F0(dummy_355_), .F1(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ), .F2(dummy_374_), .F3(\coefcal1_divide_inst1_u110_XORCI_9|SUM_net ) );
      defparam ii3436.CONFIG_DATA = 16'hEFE0;
      defparam ii3436.PLACE_LOCATION = "NONE";
      defparam ii3436.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3437 ( .DX(nn3437), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2372_), .F3(dummy_abc_2373_) );
      defparam ii3437.CONFIG_DATA = 16'h9999;
      defparam ii3437.PLACE_LOCATION = "NONE";
      defparam ii3437.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3438 ( .DX(nn3438), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_374_) );
      defparam ii3438.CONFIG_DATA = 16'hA569;
      defparam ii3438.PLACE_LOCATION = "NONE";
      defparam ii3438.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3439 ( .DX(nn3439), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_374_), .F2(nn3392), .F3(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ) );
      defparam ii3439.CONFIG_DATA = 16'hA695;
      defparam ii3439.PLACE_LOCATION = "NONE";
      defparam ii3439.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3440 ( .DX(nn3440), .F0(nn3393), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_2|SUM_net ), .F3(dummy_abc_2374_) );
      defparam ii3440.CONFIG_DATA = 16'hB8B8;
      defparam ii3440.PLACE_LOCATION = "NONE";
      defparam ii3440.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3441 ( .DX(nn3441), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3440), .F2(dummy_abc_2375_), .F3(dummy_abc_2376_) );
      defparam ii3441.CONFIG_DATA = 16'h9999;
      defparam ii3441.PLACE_LOCATION = "NONE";
      defparam ii3441.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3442 ( .DX(nn3442), .F0(nn3394), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_3|SUM_net ), .F3(dummy_abc_2377_) );
      defparam ii3442.CONFIG_DATA = 16'hB8B8;
      defparam ii3442.PLACE_LOCATION = "NONE";
      defparam ii3442.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3443 ( .DX(nn3443), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3442), .F2(dummy_abc_2378_), .F3(dummy_abc_2379_) );
      defparam ii3443.CONFIG_DATA = 16'h9999;
      defparam ii3443.PLACE_LOCATION = "NONE";
      defparam ii3443.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3444 ( .DX(nn3444), .F0(nn3395), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_4|SUM_net ), .F3(dummy_abc_2380_) );
      defparam ii3444.CONFIG_DATA = 16'hB8B8;
      defparam ii3444.PLACE_LOCATION = "NONE";
      defparam ii3444.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3445 ( .DX(nn3445), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3444), .F2(dummy_abc_2381_), .F3(dummy_abc_2382_) );
      defparam ii3445.CONFIG_DATA = 16'h9999;
      defparam ii3445.PLACE_LOCATION = "NONE";
      defparam ii3445.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3446 ( .DX(nn3446), .F0(nn3396), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_5|SUM_net ), .F3(dummy_abc_2383_) );
      defparam ii3446.CONFIG_DATA = 16'hB8B8;
      defparam ii3446.PLACE_LOCATION = "NONE";
      defparam ii3446.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3447 ( .DX(nn3447), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3446), .F2(dummy_abc_2384_), .F3(dummy_abc_2385_) );
      defparam ii3447.CONFIG_DATA = 16'h9999;
      defparam ii3447.PLACE_LOCATION = "NONE";
      defparam ii3447.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3448 ( .DX(nn3448), .F0(nn3397), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_6|SUM_net ), .F3(dummy_abc_2386_) );
      defparam ii3448.CONFIG_DATA = 16'hB8B8;
      defparam ii3448.PLACE_LOCATION = "NONE";
      defparam ii3448.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3449 ( .DX(nn3449), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3448), .F2(dummy_abc_2387_), .F3(dummy_abc_2388_) );
      defparam ii3449.CONFIG_DATA = 16'h9999;
      defparam ii3449.PLACE_LOCATION = "NONE";
      defparam ii3449.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3450 ( .DX(nn3450), .F0(nn3398), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_7|SUM_net ), .F3(dummy_abc_2389_) );
      defparam ii3450.CONFIG_DATA = 16'hB8B8;
      defparam ii3450.PLACE_LOCATION = "NONE";
      defparam ii3450.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3451 ( .DX(nn3451), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3450), .F2(dummy_abc_2390_), .F3(dummy_abc_2391_) );
      defparam ii3451.CONFIG_DATA = 16'h9999;
      defparam ii3451.PLACE_LOCATION = "NONE";
      defparam ii3451.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3452 ( .DX(nn3452), .F0(nn3399), .F1(dummy_374_), .F2(\coefcal1_divide_inst1_u110_XORCI_8|SUM_net ), .F3(dummy_abc_2392_) );
      defparam ii3452.CONFIG_DATA = 16'hB8B8;
      defparam ii3452.PLACE_LOCATION = "NONE";
      defparam ii3452.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3453 ( .DX(nn3453), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3452), .F2(dummy_abc_2393_), .F3(dummy_abc_2394_) );
      defparam ii3453.CONFIG_DATA = 16'h9999;
      defparam ii3453.PLACE_LOCATION = "NONE";
      defparam ii3453.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3454 ( .DX(nn3454), .F0(dummy_355_), .F1(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ), .F2(dummy_abc_2395_), .F3(dummy_abc_2396_) );
      defparam ii3454.CONFIG_DATA = 16'h1111;
      defparam ii3454.PLACE_LOCATION = "NONE";
      defparam ii3454.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3455 ( .DX(nn3455), .F0(nn3271), .F1(nn3454), .F2(dummy_374_), .F3(\coefcal1_divide_inst1_u110_XORCI_9|SUM_net ) );
      defparam ii3455.CONFIG_DATA = 16'h2A20;
      defparam ii3455.PLACE_LOCATION = "NONE";
      defparam ii3455.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3456 ( .DX(nn3456), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3455), .F2(dummy_abc_2397_), .F3(dummy_abc_2398_) );
      defparam ii3456.CONFIG_DATA = 16'h9999;
      defparam ii3456.PLACE_LOCATION = "NONE";
      defparam ii3456.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3457 ( .DX(nn3457), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2399_), .F2(dummy_abc_2400_), .F3(dummy_abc_2401_) );
      defparam ii3457.CONFIG_DATA = 16'h5555;
      defparam ii3457.PLACE_LOCATION = "NONE";
      defparam ii3457.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3458 ( .DX(nn3458), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2402_), .F2(dummy_abc_2403_), .F3(dummy_abc_2404_) );
      defparam ii3458.CONFIG_DATA = 16'h5555;
      defparam ii3458.PLACE_LOCATION = "NONE";
      defparam ii3458.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3459 ( .DX(nn3459), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2405_), .F2(dummy_abc_2406_), .F3(dummy_abc_2407_) );
      defparam ii3459.CONFIG_DATA = 16'h5555;
      defparam ii3459.PLACE_LOCATION = "NONE";
      defparam ii3459.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3460 ( .DX(nn3460), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2408_), .F2(dummy_abc_2409_), .F3(dummy_abc_2410_) );
      defparam ii3460.CONFIG_DATA = 16'h5555;
      defparam ii3460.PLACE_LOCATION = "NONE";
      defparam ii3460.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3461 ( .DX(nn3461), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2411_), .F2(dummy_abc_2412_), .F3(dummy_abc_2413_) );
      defparam ii3461.CONFIG_DATA = 16'h5555;
      defparam ii3461.PLACE_LOCATION = "NONE";
      defparam ii3461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3462 ( .DX(nn3462), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2414_), .F2(dummy_abc_2415_), .F3(dummy_abc_2416_) );
      defparam ii3462.CONFIG_DATA = 16'h5555;
      defparam ii3462.PLACE_LOCATION = "NONE";
      defparam ii3462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3463 ( .DX(nn3463), .F0(dummy_abc_2417_), .F1(dummy_abc_2418_), .F2(dummy_abc_2419_), .F3(dummy_abc_2420_) );
      defparam ii3463.CONFIG_DATA = 16'hFFFF;
      defparam ii3463.PLACE_LOCATION = "NONE";
      defparam ii3463.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_33_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_393_ ), 
        .DX( {nn3463, nn3462, nn3461, nn3460, nn3459, nn3458, nn3457, nn3456, 
              nn3453, nn3451, nn3449, nn3447, nn3445, nn3443, nn3441, nn3439, 
              nn3438, nn3437} ), 
        .SUM( {\coefcal1_divide_inst1_u138_XORCI_17|SUM_net , dummy_394_, 
              dummy_395_, dummy_396_, dummy_397_, dummy_398_, dummy_399_, dummy_400_, 
              dummy_401_, dummy_402_, dummy_403_, dummy_404_, dummy_405_, dummy_406_, 
              dummy_407_, dummy_408_, dummy_409_, dummy_410_} )
      );
    CS_LUT4_PRIM ii3484 ( .DX(nn3484), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_374_), .F3(dummy_abc_2421_) );
      defparam ii3484.CONFIG_DATA = 16'hA6A6;
      defparam ii3484.PLACE_LOCATION = "NONE";
      defparam ii3484.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3485 ( .DX(nn3485), .F0(dummy_374_), .F1(nn3392), .F2(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ), .F3(dummy_abc_2422_) );
      defparam ii3485.CONFIG_DATA = 16'hD8D8;
      defparam ii3485.PLACE_LOCATION = "NONE";
      defparam ii3485.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3486 ( .DX(nn3486), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2423_), .F3(dummy_abc_2424_) );
      defparam ii3486.CONFIG_DATA = 16'h9999;
      defparam ii3486.PLACE_LOCATION = "NONE";
      defparam ii3486.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3487 ( .DX(nn3487), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_374_) );
      defparam ii3487.CONFIG_DATA = 16'hA569;
      defparam ii3487.PLACE_LOCATION = "NONE";
      defparam ii3487.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3488 ( .DX(nn3488), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_374_), .F2(nn3392), .F3(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ) );
      defparam ii3488.CONFIG_DATA = 16'hA695;
      defparam ii3488.PLACE_LOCATION = "NONE";
      defparam ii3488.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3489 ( .DX(nn3489), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3440), .F2(dummy_abc_2425_), .F3(dummy_abc_2426_) );
      defparam ii3489.CONFIG_DATA = 16'h9999;
      defparam ii3489.PLACE_LOCATION = "NONE";
      defparam ii3489.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3490 ( .DX(nn3490), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3442), .F2(dummy_abc_2427_), .F3(dummy_abc_2428_) );
      defparam ii3490.CONFIG_DATA = 16'h9999;
      defparam ii3490.PLACE_LOCATION = "NONE";
      defparam ii3490.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3491 ( .DX(nn3491), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3444), .F2(dummy_abc_2429_), .F3(dummy_abc_2430_) );
      defparam ii3491.CONFIG_DATA = 16'h9999;
      defparam ii3491.PLACE_LOCATION = "NONE";
      defparam ii3491.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3492 ( .DX(nn3492), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3446), .F2(dummy_abc_2431_), .F3(dummy_abc_2432_) );
      defparam ii3492.CONFIG_DATA = 16'h9999;
      defparam ii3492.PLACE_LOCATION = "NONE";
      defparam ii3492.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3493 ( .DX(nn3493), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3448), .F2(dummy_abc_2433_), .F3(dummy_abc_2434_) );
      defparam ii3493.CONFIG_DATA = 16'h9999;
      defparam ii3493.PLACE_LOCATION = "NONE";
      defparam ii3493.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3494 ( .DX(nn3494), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3450), .F2(dummy_abc_2435_), .F3(dummy_abc_2436_) );
      defparam ii3494.CONFIG_DATA = 16'h9999;
      defparam ii3494.PLACE_LOCATION = "NONE";
      defparam ii3494.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3495 ( .DX(nn3495), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3452), .F2(dummy_abc_2437_), .F3(dummy_abc_2438_) );
      defparam ii3495.CONFIG_DATA = 16'h9999;
      defparam ii3495.PLACE_LOCATION = "NONE";
      defparam ii3495.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3496 ( .DX(nn3496), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3455), .F2(dummy_abc_2439_), .F3(dummy_abc_2440_) );
      defparam ii3496.CONFIG_DATA = 16'h9999;
      defparam ii3496.PLACE_LOCATION = "NONE";
      defparam ii3496.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3497 ( .DX(nn3497), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2441_), .F2(dummy_abc_2442_), .F3(dummy_abc_2443_) );
      defparam ii3497.CONFIG_DATA = 16'h5555;
      defparam ii3497.PLACE_LOCATION = "NONE";
      defparam ii3497.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3498 ( .DX(nn3498), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2444_), .F2(dummy_abc_2445_), .F3(dummy_abc_2446_) );
      defparam ii3498.CONFIG_DATA = 16'h5555;
      defparam ii3498.PLACE_LOCATION = "NONE";
      defparam ii3498.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3499 ( .DX(nn3499), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2447_), .F2(dummy_abc_2448_), .F3(dummy_abc_2449_) );
      defparam ii3499.CONFIG_DATA = 16'h5555;
      defparam ii3499.PLACE_LOCATION = "NONE";
      defparam ii3499.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3500 ( .DX(nn3500), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2450_), .F2(dummy_abc_2451_), .F3(dummy_abc_2452_) );
      defparam ii3500.CONFIG_DATA = 16'h5555;
      defparam ii3500.PLACE_LOCATION = "NONE";
      defparam ii3500.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3501 ( .DX(nn3501), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2453_), .F2(dummy_abc_2454_), .F3(dummy_abc_2455_) );
      defparam ii3501.CONFIG_DATA = 16'h5555;
      defparam ii3501.PLACE_LOCATION = "NONE";
      defparam ii3501.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3502 ( .DX(nn3502), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2456_), .F2(dummy_abc_2457_), .F3(dummy_abc_2458_) );
      defparam ii3502.CONFIG_DATA = 16'h5555;
      defparam ii3502.PLACE_LOCATION = "NONE";
      defparam ii3502.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_18_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn3455, nn3452, nn3450, nn3448, nn3446, nn3444, nn3442, 
              nn3440, nn3485, nn3484, \coefcal1_xDividend__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_156_ ), 
        .DX( {nn3502, nn3501, nn3500, nn3499, nn3498, nn3497, nn3496, nn3495, 
              nn3494, nn3493, nn3492, nn3491, nn3490, nn3489, nn3488, nn3487, 
              nn3486} ), 
        .SUM( {dummy_157_, \coefcal1_divide_inst1_u111_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_14|SUM_net , \coefcal1_divide_inst1_u111_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_12|SUM_net , \coefcal1_divide_inst1_u111_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_10|SUM_net , \coefcal1_divide_inst1_u111_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_8|SUM_net , \coefcal1_divide_inst1_u111_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_6|SUM_net , \coefcal1_divide_inst1_u111_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_4|SUM_net , \coefcal1_divide_inst1_u111_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_2|SUM_net , \coefcal1_divide_inst1_u111_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3522 ( .DX(nn3522), .F0(nn3271), .F1(nn3436), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_10|SUM_net ) );
      defparam ii3522.CONFIG_DATA = 16'h8A80;
      defparam ii3522.PLACE_LOCATION = "NONE";
      defparam ii3522.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3523 ( .DX(nn3523), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2459_), .F3(dummy_abc_2460_) );
      defparam ii3523.CONFIG_DATA = 16'h9999;
      defparam ii3523.PLACE_LOCATION = "NONE";
      defparam ii3523.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3524 ( .DX(nn3524), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_393_) );
      defparam ii3524.CONFIG_DATA = 16'hA569;
      defparam ii3524.PLACE_LOCATION = "NONE";
      defparam ii3524.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3525 ( .DX(nn3525), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_393_), .F2(nn3484), .F3(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ) );
      defparam ii3525.CONFIG_DATA = 16'hA695;
      defparam ii3525.PLACE_LOCATION = "NONE";
      defparam ii3525.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3526 ( .DX(nn3526), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3485), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ) );
      defparam ii3526.CONFIG_DATA = 16'h9A95;
      defparam ii3526.PLACE_LOCATION = "NONE";
      defparam ii3526.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3527 ( .DX(nn3527), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3440), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ) );
      defparam ii3527.CONFIG_DATA = 16'h9A95;
      defparam ii3527.PLACE_LOCATION = "NONE";
      defparam ii3527.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3528 ( .DX(nn3528), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3442), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ) );
      defparam ii3528.CONFIG_DATA = 16'h9A95;
      defparam ii3528.PLACE_LOCATION = "NONE";
      defparam ii3528.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3529 ( .DX(nn3529), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3444), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ) );
      defparam ii3529.CONFIG_DATA = 16'h9A95;
      defparam ii3529.PLACE_LOCATION = "NONE";
      defparam ii3529.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3530 ( .DX(nn3530), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3446), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ) );
      defparam ii3530.CONFIG_DATA = 16'h9A95;
      defparam ii3530.PLACE_LOCATION = "NONE";
      defparam ii3530.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3531 ( .DX(nn3531), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3448), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ) );
      defparam ii3531.CONFIG_DATA = 16'h9A95;
      defparam ii3531.PLACE_LOCATION = "NONE";
      defparam ii3531.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3532 ( .DX(nn3532), .F0(nn3450), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_8|SUM_net ), .F3(dummy_abc_2461_) );
      defparam ii3532.CONFIG_DATA = 16'hB8B8;
      defparam ii3532.PLACE_LOCATION = "NONE";
      defparam ii3532.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3533 ( .DX(nn3533), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3532), .F2(dummy_abc_2462_), .F3(dummy_abc_2463_) );
      defparam ii3533.CONFIG_DATA = 16'h9999;
      defparam ii3533.PLACE_LOCATION = "NONE";
      defparam ii3533.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3534 ( .DX(nn3534), .F0(nn3452), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_9|SUM_net ), .F3(dummy_abc_2464_) );
      defparam ii3534.CONFIG_DATA = 16'hB8B8;
      defparam ii3534.PLACE_LOCATION = "NONE";
      defparam ii3534.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3535 ( .DX(nn3535), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3534), .F2(dummy_abc_2465_), .F3(dummy_abc_2466_) );
      defparam ii3535.CONFIG_DATA = 16'h9999;
      defparam ii3535.PLACE_LOCATION = "NONE";
      defparam ii3535.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3536 ( .DX(nn3536), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3522), .F2(dummy_abc_2467_), .F3(dummy_abc_2468_) );
      defparam ii3536.CONFIG_DATA = 16'h9999;
      defparam ii3536.PLACE_LOCATION = "NONE";
      defparam ii3536.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3537 ( .DX(nn3537), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2469_), .F2(dummy_abc_2470_), .F3(dummy_abc_2471_) );
      defparam ii3537.CONFIG_DATA = 16'h5555;
      defparam ii3537.PLACE_LOCATION = "NONE";
      defparam ii3537.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3538 ( .DX(nn3538), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2472_), .F2(dummy_abc_2473_), .F3(dummy_abc_2474_) );
      defparam ii3538.CONFIG_DATA = 16'h5555;
      defparam ii3538.PLACE_LOCATION = "NONE";
      defparam ii3538.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3539 ( .DX(nn3539), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2475_), .F2(dummy_abc_2476_), .F3(dummy_abc_2477_) );
      defparam ii3539.CONFIG_DATA = 16'h5555;
      defparam ii3539.PLACE_LOCATION = "NONE";
      defparam ii3539.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3540 ( .DX(nn3540), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2478_), .F2(dummy_abc_2479_), .F3(dummy_abc_2480_) );
      defparam ii3540.CONFIG_DATA = 16'h5555;
      defparam ii3540.PLACE_LOCATION = "NONE";
      defparam ii3540.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3541 ( .DX(nn3541), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2481_), .F2(dummy_abc_2482_), .F3(dummy_abc_2483_) );
      defparam ii3541.CONFIG_DATA = 16'h5555;
      defparam ii3541.PLACE_LOCATION = "NONE";
      defparam ii3541.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3542 ( .DX(nn3542), .F0(dummy_abc_2484_), .F1(dummy_abc_2485_), .F2(dummy_abc_2486_), .F3(dummy_abc_2487_) );
      defparam ii3542.CONFIG_DATA = 16'hFFFF;
      defparam ii3542.PLACE_LOCATION = "NONE";
      defparam ii3542.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_34_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_412_ ), 
        .DX( {nn3542, nn3541, nn3540, nn3539, nn3538, nn3537, nn3536, nn3535, 
              nn3533, nn3531, nn3530, nn3529, nn3528, nn3527, nn3526, nn3525, 
              nn3524, nn3523} ), 
        .SUM( {\coefcal1_divide_inst1_u140_XORCI_17|SUM_net , dummy_413_, 
              dummy_414_, dummy_415_, dummy_416_, dummy_417_, dummy_418_, dummy_419_, 
              dummy_420_, dummy_421_, dummy_422_, dummy_423_, dummy_424_, dummy_425_, 
              dummy_426_, dummy_427_, dummy_428_, dummy_429_} )
      );
    CS_LUT4_PRIM ii3563 ( .DX(nn3563), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2488_), .F3(dummy_abc_2489_) );
      defparam ii3563.CONFIG_DATA = 16'h9999;
      defparam ii3563.PLACE_LOCATION = "NONE";
      defparam ii3563.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3564 ( .DX(nn3564), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_412_) );
      defparam ii3564.CONFIG_DATA = 16'hA569;
      defparam ii3564.PLACE_LOCATION = "NONE";
      defparam ii3564.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3565 ( .DX(nn3565), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_393_), .F3(dummy_abc_2490_) );
      defparam ii3565.CONFIG_DATA = 16'hA6A6;
      defparam ii3565.PLACE_LOCATION = "NONE";
      defparam ii3565.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3566 ( .DX(nn3566), .F0(dummy_393_), .F1(nn3484), .F2(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ), .F3(dummy_abc_2491_) );
      defparam ii3566.CONFIG_DATA = 16'hD8D8;
      defparam ii3566.PLACE_LOCATION = "NONE";
      defparam ii3566.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3567 ( .DX(nn3567), .F0(nn3485), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ), .F3(dummy_abc_2492_) );
      defparam ii3567.CONFIG_DATA = 16'hB8B8;
      defparam ii3567.PLACE_LOCATION = "NONE";
      defparam ii3567.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3568 ( .DX(nn3568), .F0(nn3440), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ), .F3(dummy_abc_2493_) );
      defparam ii3568.CONFIG_DATA = 16'hB8B8;
      defparam ii3568.PLACE_LOCATION = "NONE";
      defparam ii3568.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3569 ( .DX(nn3569), .F0(nn3442), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ), .F3(dummy_abc_2494_) );
      defparam ii3569.CONFIG_DATA = 16'hB8B8;
      defparam ii3569.PLACE_LOCATION = "NONE";
      defparam ii3569.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3570 ( .DX(nn3570), .F0(nn3444), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ), .F3(dummy_abc_2495_) );
      defparam ii3570.CONFIG_DATA = 16'hB8B8;
      defparam ii3570.PLACE_LOCATION = "NONE";
      defparam ii3570.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3571 ( .DX(nn3571), .F0(nn3446), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ), .F3(dummy_abc_2496_) );
      defparam ii3571.CONFIG_DATA = 16'hB8B8;
      defparam ii3571.PLACE_LOCATION = "NONE";
      defparam ii3571.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3572 ( .DX(nn3572), .F0(nn3448), .F1(dummy_393_), .F2(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ), .F3(dummy_abc_2497_) );
      defparam ii3572.CONFIG_DATA = 16'hB8B8;
      defparam ii3572.PLACE_LOCATION = "NONE";
      defparam ii3572.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3573 ( .DX(nn3573), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2498_), .F3(dummy_abc_2499_) );
      defparam ii3573.CONFIG_DATA = 16'h9999;
      defparam ii3573.PLACE_LOCATION = "NONE";
      defparam ii3573.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3574 ( .DX(nn3574), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_393_) );
      defparam ii3574.CONFIG_DATA = 16'hA569;
      defparam ii3574.PLACE_LOCATION = "NONE";
      defparam ii3574.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3575 ( .DX(nn3575), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_393_), .F2(nn3484), .F3(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ) );
      defparam ii3575.CONFIG_DATA = 16'hA695;
      defparam ii3575.PLACE_LOCATION = "NONE";
      defparam ii3575.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3576 ( .DX(nn3576), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3485), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ) );
      defparam ii3576.CONFIG_DATA = 16'h9A95;
      defparam ii3576.PLACE_LOCATION = "NONE";
      defparam ii3576.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3577 ( .DX(nn3577), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3440), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ) );
      defparam ii3577.CONFIG_DATA = 16'h9A95;
      defparam ii3577.PLACE_LOCATION = "NONE";
      defparam ii3577.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3578 ( .DX(nn3578), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3442), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ) );
      defparam ii3578.CONFIG_DATA = 16'h9A95;
      defparam ii3578.PLACE_LOCATION = "NONE";
      defparam ii3578.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3579 ( .DX(nn3579), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3444), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ) );
      defparam ii3579.CONFIG_DATA = 16'h9A95;
      defparam ii3579.PLACE_LOCATION = "NONE";
      defparam ii3579.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3580 ( .DX(nn3580), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3446), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ) );
      defparam ii3580.CONFIG_DATA = 16'h9A95;
      defparam ii3580.PLACE_LOCATION = "NONE";
      defparam ii3580.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3581 ( .DX(nn3581), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3448), .F2(dummy_393_), .F3(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ) );
      defparam ii3581.CONFIG_DATA = 16'h9A95;
      defparam ii3581.PLACE_LOCATION = "NONE";
      defparam ii3581.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3582 ( .DX(nn3582), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3532), .F2(dummy_abc_2500_), .F3(dummy_abc_2501_) );
      defparam ii3582.CONFIG_DATA = 16'h9999;
      defparam ii3582.PLACE_LOCATION = "NONE";
      defparam ii3582.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3583 ( .DX(nn3583), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3534), .F2(dummy_abc_2502_), .F3(dummy_abc_2503_) );
      defparam ii3583.CONFIG_DATA = 16'h9999;
      defparam ii3583.PLACE_LOCATION = "NONE";
      defparam ii3583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3584 ( .DX(nn3584), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3522), .F2(dummy_abc_2504_), .F3(dummy_abc_2505_) );
      defparam ii3584.CONFIG_DATA = 16'h9999;
      defparam ii3584.PLACE_LOCATION = "NONE";
      defparam ii3584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3585 ( .DX(nn3585), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2506_), .F2(dummy_abc_2507_), .F3(dummy_abc_2508_) );
      defparam ii3585.CONFIG_DATA = 16'h5555;
      defparam ii3585.PLACE_LOCATION = "NONE";
      defparam ii3585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3586 ( .DX(nn3586), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2509_), .F2(dummy_abc_2510_), .F3(dummy_abc_2511_) );
      defparam ii3586.CONFIG_DATA = 16'h5555;
      defparam ii3586.PLACE_LOCATION = "NONE";
      defparam ii3586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3587 ( .DX(nn3587), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2512_), .F2(dummy_abc_2513_), .F3(dummy_abc_2514_) );
      defparam ii3587.CONFIG_DATA = 16'h5555;
      defparam ii3587.PLACE_LOCATION = "NONE";
      defparam ii3587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3588 ( .DX(nn3588), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2515_), .F2(dummy_abc_2516_), .F3(dummy_abc_2517_) );
      defparam ii3588.CONFIG_DATA = 16'h5555;
      defparam ii3588.PLACE_LOCATION = "NONE";
      defparam ii3588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3589 ( .DX(nn3589), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2518_), .F2(dummy_abc_2519_), .F3(dummy_abc_2520_) );
      defparam ii3589.CONFIG_DATA = 16'h5555;
      defparam ii3589.PLACE_LOCATION = "NONE";
      defparam ii3589.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_19_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3522, 
              nn3534, nn3532, nn3572, nn3571, nn3570, nn3569, nn3568, nn3567, 
              nn3566, nn3565, \coefcal1_xDividend__reg[5]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_158_ ), 
        .DX( {nn3589, nn3588, nn3587, nn3586, nn3585, nn3584, nn3583, nn3582, 
              nn3581, nn3580, nn3579, nn3578, nn3577, nn3576, nn3575, nn3574, 
              nn3573} ), 
        .SUM( {dummy_159_, \coefcal1_divide_inst1_u112_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_14|SUM_net , \coefcal1_divide_inst1_u112_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_12|SUM_net , \coefcal1_divide_inst1_u112_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_10|SUM_net , \coefcal1_divide_inst1_u112_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_8|SUM_net , \coefcal1_divide_inst1_u112_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_6|SUM_net , \coefcal1_divide_inst1_u112_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_4|SUM_net , \coefcal1_divide_inst1_u112_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_2|SUM_net , \coefcal1_divide_inst1_u112_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3609 ( .DX(nn3609), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_412_), .F2(nn3565), .F3(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ) );
      defparam ii3609.CONFIG_DATA = 16'hA695;
      defparam ii3609.PLACE_LOCATION = "NONE";
      defparam ii3609.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3610 ( .DX(nn3610), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3566), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ) );
      defparam ii3610.CONFIG_DATA = 16'h9A95;
      defparam ii3610.PLACE_LOCATION = "NONE";
      defparam ii3610.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3611 ( .DX(nn3611), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3567), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ) );
      defparam ii3611.CONFIG_DATA = 16'h9A95;
      defparam ii3611.PLACE_LOCATION = "NONE";
      defparam ii3611.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3612 ( .DX(nn3612), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3568), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ) );
      defparam ii3612.CONFIG_DATA = 16'h9A95;
      defparam ii3612.PLACE_LOCATION = "NONE";
      defparam ii3612.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3613 ( .DX(nn3613), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3569), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ) );
      defparam ii3613.CONFIG_DATA = 16'h9A95;
      defparam ii3613.PLACE_LOCATION = "NONE";
      defparam ii3613.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3614 ( .DX(nn3614), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3570), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ) );
      defparam ii3614.CONFIG_DATA = 16'h9A95;
      defparam ii3614.PLACE_LOCATION = "NONE";
      defparam ii3614.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3615 ( .DX(nn3615), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3571), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ) );
      defparam ii3615.CONFIG_DATA = 16'h9A95;
      defparam ii3615.PLACE_LOCATION = "NONE";
      defparam ii3615.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3616 ( .DX(nn3616), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3572), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ) );
      defparam ii3616.CONFIG_DATA = 16'h9A95;
      defparam ii3616.PLACE_LOCATION = "NONE";
      defparam ii3616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3617 ( .DX(nn3617), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3532), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ) );
      defparam ii3617.CONFIG_DATA = 16'h9A95;
      defparam ii3617.PLACE_LOCATION = "NONE";
      defparam ii3617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3618 ( .DX(nn3618), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3534), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ) );
      defparam ii3618.CONFIG_DATA = 16'h9A95;
      defparam ii3618.PLACE_LOCATION = "NONE";
      defparam ii3618.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3619 ( .DX(nn3619), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3522), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_11|SUM_net ) );
      defparam ii3619.CONFIG_DATA = 16'h9A95;
      defparam ii3619.PLACE_LOCATION = "NONE";
      defparam ii3619.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3620 ( .DX(nn3620), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2521_), .F2(dummy_abc_2522_), .F3(dummy_abc_2523_) );
      defparam ii3620.CONFIG_DATA = 16'h5555;
      defparam ii3620.PLACE_LOCATION = "NONE";
      defparam ii3620.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3621 ( .DX(nn3621), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2524_), .F2(dummy_abc_2525_), .F3(dummy_abc_2526_) );
      defparam ii3621.CONFIG_DATA = 16'h5555;
      defparam ii3621.PLACE_LOCATION = "NONE";
      defparam ii3621.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3622 ( .DX(nn3622), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2527_), .F2(dummy_abc_2528_), .F3(dummy_abc_2529_) );
      defparam ii3622.CONFIG_DATA = 16'h5555;
      defparam ii3622.PLACE_LOCATION = "NONE";
      defparam ii3622.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3623 ( .DX(nn3623), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2530_), .F2(dummy_abc_2531_), .F3(dummy_abc_2532_) );
      defparam ii3623.CONFIG_DATA = 16'h5555;
      defparam ii3623.PLACE_LOCATION = "NONE";
      defparam ii3623.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3624 ( .DX(nn3624), .F0(dummy_abc_2533_), .F1(dummy_abc_2534_), .F2(dummy_abc_2535_), .F3(dummy_abc_2536_) );
      defparam ii3624.CONFIG_DATA = 16'hFFFF;
      defparam ii3624.PLACE_LOCATION = "NONE";
      defparam ii3624.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_35_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_431_ ), 
        .DX( {nn3624, nn3623, nn3622, nn3621, nn3620, nn3619, nn3618, nn3617, 
              nn3616, nn3615, nn3614, nn3613, nn3612, nn3611, nn3610, nn3609, 
              nn3564, nn3563} ), 
        .SUM( {\coefcal1_divide_inst1_u142_XORCI_17|SUM_net , dummy_432_, 
              dummy_433_, dummy_434_, dummy_435_, dummy_436_, dummy_437_, dummy_438_, 
              dummy_439_, dummy_440_, dummy_441_, dummy_442_, dummy_443_, dummy_444_, 
              dummy_445_, dummy_446_, dummy_447_, dummy_448_} )
      );
    CS_LUT4_PRIM ii3645 ( .DX(nn3645), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_412_), .F3(dummy_abc_2537_) );
      defparam ii3645.CONFIG_DATA = 16'hA6A6;
      defparam ii3645.PLACE_LOCATION = "NONE";
      defparam ii3645.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3646 ( .DX(nn3646), .F0(dummy_412_), .F1(nn3565), .F2(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ), .F3(dummy_abc_2538_) );
      defparam ii3646.CONFIG_DATA = 16'hD8D8;
      defparam ii3646.PLACE_LOCATION = "NONE";
      defparam ii3646.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3647 ( .DX(nn3647), .F0(nn3566), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ), .F3(dummy_abc_2539_) );
      defparam ii3647.CONFIG_DATA = 16'hB8B8;
      defparam ii3647.PLACE_LOCATION = "NONE";
      defparam ii3647.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3648 ( .DX(nn3648), .F0(nn3567), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ), .F3(dummy_abc_2540_) );
      defparam ii3648.CONFIG_DATA = 16'hB8B8;
      defparam ii3648.PLACE_LOCATION = "NONE";
      defparam ii3648.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3649 ( .DX(nn3649), .F0(nn3568), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ), .F3(dummy_abc_2541_) );
      defparam ii3649.CONFIG_DATA = 16'hB8B8;
      defparam ii3649.PLACE_LOCATION = "NONE";
      defparam ii3649.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3650 ( .DX(nn3650), .F0(nn3569), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ), .F3(dummy_abc_2542_) );
      defparam ii3650.CONFIG_DATA = 16'hB8B8;
      defparam ii3650.PLACE_LOCATION = "NONE";
      defparam ii3650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3651 ( .DX(nn3651), .F0(nn3570), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ), .F3(dummy_abc_2543_) );
      defparam ii3651.CONFIG_DATA = 16'hB8B8;
      defparam ii3651.PLACE_LOCATION = "NONE";
      defparam ii3651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3652 ( .DX(nn3652), .F0(nn3571), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ), .F3(dummy_abc_2544_) );
      defparam ii3652.CONFIG_DATA = 16'hB8B8;
      defparam ii3652.PLACE_LOCATION = "NONE";
      defparam ii3652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3653 ( .DX(nn3653), .F0(nn3572), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ), .F3(dummy_abc_2545_) );
      defparam ii3653.CONFIG_DATA = 16'hB8B8;
      defparam ii3653.PLACE_LOCATION = "NONE";
      defparam ii3653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3654 ( .DX(nn3654), .F0(nn3532), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ), .F3(dummy_abc_2546_) );
      defparam ii3654.CONFIG_DATA = 16'hB8B8;
      defparam ii3654.PLACE_LOCATION = "NONE";
      defparam ii3654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3655 ( .DX(nn3655), .F0(nn3534), .F1(dummy_412_), .F2(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ), .F3(dummy_abc_2547_) );
      defparam ii3655.CONFIG_DATA = 16'hB8B8;
      defparam ii3655.PLACE_LOCATION = "NONE";
      defparam ii3655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3656 ( .DX(nn3656), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2548_), .F3(dummy_abc_2549_) );
      defparam ii3656.CONFIG_DATA = 16'h9999;
      defparam ii3656.PLACE_LOCATION = "NONE";
      defparam ii3656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3657 ( .DX(nn3657), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_412_) );
      defparam ii3657.CONFIG_DATA = 16'hA569;
      defparam ii3657.PLACE_LOCATION = "NONE";
      defparam ii3657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3658 ( .DX(nn3658), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_412_), .F2(nn3565), .F3(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ) );
      defparam ii3658.CONFIG_DATA = 16'hA695;
      defparam ii3658.PLACE_LOCATION = "NONE";
      defparam ii3658.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3659 ( .DX(nn3659), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3566), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ) );
      defparam ii3659.CONFIG_DATA = 16'h9A95;
      defparam ii3659.PLACE_LOCATION = "NONE";
      defparam ii3659.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3660 ( .DX(nn3660), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3567), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ) );
      defparam ii3660.CONFIG_DATA = 16'h9A95;
      defparam ii3660.PLACE_LOCATION = "NONE";
      defparam ii3660.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3661 ( .DX(nn3661), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3568), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ) );
      defparam ii3661.CONFIG_DATA = 16'h9A95;
      defparam ii3661.PLACE_LOCATION = "NONE";
      defparam ii3661.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3662 ( .DX(nn3662), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3569), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ) );
      defparam ii3662.CONFIG_DATA = 16'h9A95;
      defparam ii3662.PLACE_LOCATION = "NONE";
      defparam ii3662.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3663 ( .DX(nn3663), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3570), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ) );
      defparam ii3663.CONFIG_DATA = 16'h9A95;
      defparam ii3663.PLACE_LOCATION = "NONE";
      defparam ii3663.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3664 ( .DX(nn3664), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3571), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ) );
      defparam ii3664.CONFIG_DATA = 16'h9A95;
      defparam ii3664.PLACE_LOCATION = "NONE";
      defparam ii3664.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3665 ( .DX(nn3665), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3572), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ) );
      defparam ii3665.CONFIG_DATA = 16'h9A95;
      defparam ii3665.PLACE_LOCATION = "NONE";
      defparam ii3665.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3666 ( .DX(nn3666), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3532), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ) );
      defparam ii3666.CONFIG_DATA = 16'h9A95;
      defparam ii3666.PLACE_LOCATION = "NONE";
      defparam ii3666.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3667 ( .DX(nn3667), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3534), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ) );
      defparam ii3667.CONFIG_DATA = 16'h9A95;
      defparam ii3667.PLACE_LOCATION = "NONE";
      defparam ii3667.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3668 ( .DX(nn3668), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3522), .F2(dummy_412_), .F3(\coefcal1_divide_inst1_u112_XORCI_11|SUM_net ) );
      defparam ii3668.CONFIG_DATA = 16'h9A95;
      defparam ii3668.PLACE_LOCATION = "NONE";
      defparam ii3668.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3669 ( .DX(nn3669), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2550_), .F2(dummy_abc_2551_), .F3(dummy_abc_2552_) );
      defparam ii3669.CONFIG_DATA = 16'h5555;
      defparam ii3669.PLACE_LOCATION = "NONE";
      defparam ii3669.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3670 ( .DX(nn3670), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2553_), .F2(dummy_abc_2554_), .F3(dummy_abc_2555_) );
      defparam ii3670.CONFIG_DATA = 16'h5555;
      defparam ii3670.PLACE_LOCATION = "NONE";
      defparam ii3670.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3671 ( .DX(nn3671), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2556_), .F2(dummy_abc_2557_), .F3(dummy_abc_2558_) );
      defparam ii3671.CONFIG_DATA = 16'h5555;
      defparam ii3671.PLACE_LOCATION = "NONE";
      defparam ii3671.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3672 ( .DX(nn3672), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2559_), .F2(dummy_abc_2560_), .F3(dummy_abc_2561_) );
      defparam ii3672.CONFIG_DATA = 16'h5555;
      defparam ii3672.PLACE_LOCATION = "NONE";
      defparam ii3672.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_20_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3655, 
              nn3654, nn3653, nn3652, nn3651, nn3650, nn3649, nn3648, nn3647, 
              nn3646, nn3645, \coefcal1_xDividend__reg[4]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_160_ ), 
        .DX( {nn3672, nn3671, nn3670, nn3669, nn3668, nn3667, nn3666, nn3665, 
              nn3664, nn3663, nn3662, nn3661, nn3660, nn3659, nn3658, nn3657, 
              nn3656} ), 
        .SUM( {dummy_161_, \coefcal1_divide_inst1_u113_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_14|SUM_net , \coefcal1_divide_inst1_u113_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_12|SUM_net , \coefcal1_divide_inst1_u113_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_10|SUM_net , \coefcal1_divide_inst1_u113_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_8|SUM_net , \coefcal1_divide_inst1_u113_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_6|SUM_net , \coefcal1_divide_inst1_u113_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_4|SUM_net , \coefcal1_divide_inst1_u113_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_2|SUM_net , \coefcal1_divide_inst1_u113_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3692 ( .DX(nn3692), .F0(nn3522), .F1(dummy_412_), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3692.CONFIG_DATA = 16'h8F80;
      defparam ii3692.PLACE_LOCATION = "NONE";
      defparam ii3692.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3693 ( .DX(nn3693), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2562_), .F3(dummy_abc_2563_) );
      defparam ii3693.CONFIG_DATA = 16'h9999;
      defparam ii3693.PLACE_LOCATION = "NONE";
      defparam ii3693.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3694 ( .DX(nn3694), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_431_) );
      defparam ii3694.CONFIG_DATA = 16'hA569;
      defparam ii3694.PLACE_LOCATION = "NONE";
      defparam ii3694.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3695 ( .DX(nn3695), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_431_), .F2(nn3645), .F3(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ) );
      defparam ii3695.CONFIG_DATA = 16'hA695;
      defparam ii3695.PLACE_LOCATION = "NONE";
      defparam ii3695.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3696 ( .DX(nn3696), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3646), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ) );
      defparam ii3696.CONFIG_DATA = 16'h9A95;
      defparam ii3696.PLACE_LOCATION = "NONE";
      defparam ii3696.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3697 ( .DX(nn3697), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3647), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ) );
      defparam ii3697.CONFIG_DATA = 16'h9A95;
      defparam ii3697.PLACE_LOCATION = "NONE";
      defparam ii3697.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3698 ( .DX(nn3698), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3648), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ) );
      defparam ii3698.CONFIG_DATA = 16'h9A95;
      defparam ii3698.PLACE_LOCATION = "NONE";
      defparam ii3698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3699 ( .DX(nn3699), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3649), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ) );
      defparam ii3699.CONFIG_DATA = 16'h9A95;
      defparam ii3699.PLACE_LOCATION = "NONE";
      defparam ii3699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3700 ( .DX(nn3700), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3650), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ) );
      defparam ii3700.CONFIG_DATA = 16'h9A95;
      defparam ii3700.PLACE_LOCATION = "NONE";
      defparam ii3700.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3701 ( .DX(nn3701), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3651), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ) );
      defparam ii3701.CONFIG_DATA = 16'h9A95;
      defparam ii3701.PLACE_LOCATION = "NONE";
      defparam ii3701.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3702 ( .DX(nn3702), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3652), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ) );
      defparam ii3702.CONFIG_DATA = 16'h9A95;
      defparam ii3702.PLACE_LOCATION = "NONE";
      defparam ii3702.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3703 ( .DX(nn3703), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3653), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ) );
      defparam ii3703.CONFIG_DATA = 16'h9A95;
      defparam ii3703.PLACE_LOCATION = "NONE";
      defparam ii3703.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3704 ( .DX(nn3704), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3654), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ) );
      defparam ii3704.CONFIG_DATA = 16'h9A95;
      defparam ii3704.PLACE_LOCATION = "NONE";
      defparam ii3704.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3705 ( .DX(nn3705), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3655), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ) );
      defparam ii3705.CONFIG_DATA = 16'h9A95;
      defparam ii3705.PLACE_LOCATION = "NONE";
      defparam ii3705.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3706 ( .DX(nn3706), .F0(nn3522), .F1(dummy_412_), .F2(dummy_abc_2564_), .F3(dummy_abc_2565_) );
      defparam ii3706.CONFIG_DATA = 16'h8888;
      defparam ii3706.PLACE_LOCATION = "NONE";
      defparam ii3706.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3707 ( .DX(nn3707), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3706), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3707.CONFIG_DATA = 16'h9095;
      defparam ii3707.PLACE_LOCATION = "NONE";
      defparam ii3707.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3708 ( .DX(nn3708), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2566_), .F2(dummy_abc_2567_), .F3(dummy_abc_2568_) );
      defparam ii3708.CONFIG_DATA = 16'h5555;
      defparam ii3708.PLACE_LOCATION = "NONE";
      defparam ii3708.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3709 ( .DX(nn3709), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2569_), .F2(dummy_abc_2570_), .F3(dummy_abc_2571_) );
      defparam ii3709.CONFIG_DATA = 16'h5555;
      defparam ii3709.PLACE_LOCATION = "NONE";
      defparam ii3709.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3710 ( .DX(nn3710), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2572_), .F2(dummy_abc_2573_), .F3(dummy_abc_2574_) );
      defparam ii3710.CONFIG_DATA = 16'h5555;
      defparam ii3710.PLACE_LOCATION = "NONE";
      defparam ii3710.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3711 ( .DX(nn3711), .F0(dummy_abc_2575_), .F1(dummy_abc_2576_), .F2(dummy_abc_2577_), .F3(dummy_abc_2578_) );
      defparam ii3711.CONFIG_DATA = 16'hFFFF;
      defparam ii3711.PLACE_LOCATION = "NONE";
      defparam ii3711.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_36_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_450_ ), 
        .DX( {nn3711, nn3710, nn3709, nn3708, nn3707, nn3705, nn3704, nn3703, 
              nn3702, nn3701, nn3700, nn3699, nn3698, nn3697, nn3696, nn3695, 
              nn3694, nn3693} ), 
        .SUM( {\coefcal1_divide_inst1_u144_XORCI_17|SUM_net , dummy_451_, 
              dummy_452_, dummy_453_, dummy_454_, dummy_455_, dummy_456_, dummy_457_, 
              dummy_458_, dummy_459_, dummy_460_, dummy_461_, dummy_462_, dummy_463_, 
              dummy_464_, dummy_465_, dummy_466_, dummy_467_} )
      );
    CS_LUT4_PRIM ii3732 ( .DX(nn3732), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_431_), .F3(dummy_abc_2579_) );
      defparam ii3732.CONFIG_DATA = 16'hA6A6;
      defparam ii3732.PLACE_LOCATION = "NONE";
      defparam ii3732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3733 ( .DX(nn3733), .F0(dummy_431_), .F1(nn3645), .F2(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ), .F3(dummy_abc_2580_) );
      defparam ii3733.CONFIG_DATA = 16'hD8D8;
      defparam ii3733.PLACE_LOCATION = "NONE";
      defparam ii3733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3734 ( .DX(nn3734), .F0(nn3646), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ), .F3(dummy_abc_2581_) );
      defparam ii3734.CONFIG_DATA = 16'hB8B8;
      defparam ii3734.PLACE_LOCATION = "NONE";
      defparam ii3734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3735 ( .DX(nn3735), .F0(nn3647), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ), .F3(dummy_abc_2582_) );
      defparam ii3735.CONFIG_DATA = 16'hB8B8;
      defparam ii3735.PLACE_LOCATION = "NONE";
      defparam ii3735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3736 ( .DX(nn3736), .F0(nn3648), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ), .F3(dummy_abc_2583_) );
      defparam ii3736.CONFIG_DATA = 16'hB8B8;
      defparam ii3736.PLACE_LOCATION = "NONE";
      defparam ii3736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3737 ( .DX(nn3737), .F0(nn3649), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ), .F3(dummy_abc_2584_) );
      defparam ii3737.CONFIG_DATA = 16'hB8B8;
      defparam ii3737.PLACE_LOCATION = "NONE";
      defparam ii3737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3738 ( .DX(nn3738), .F0(nn3650), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ), .F3(dummy_abc_2585_) );
      defparam ii3738.CONFIG_DATA = 16'hB8B8;
      defparam ii3738.PLACE_LOCATION = "NONE";
      defparam ii3738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3739 ( .DX(nn3739), .F0(nn3651), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ), .F3(dummy_abc_2586_) );
      defparam ii3739.CONFIG_DATA = 16'hB8B8;
      defparam ii3739.PLACE_LOCATION = "NONE";
      defparam ii3739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3740 ( .DX(nn3740), .F0(nn3652), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ), .F3(dummy_abc_2587_) );
      defparam ii3740.CONFIG_DATA = 16'hB8B8;
      defparam ii3740.PLACE_LOCATION = "NONE";
      defparam ii3740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3741 ( .DX(nn3741), .F0(nn3653), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ), .F3(dummy_abc_2588_) );
      defparam ii3741.CONFIG_DATA = 16'hB8B8;
      defparam ii3741.PLACE_LOCATION = "NONE";
      defparam ii3741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3742 ( .DX(nn3742), .F0(nn3654), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ), .F3(dummy_abc_2589_) );
      defparam ii3742.CONFIG_DATA = 16'hB8B8;
      defparam ii3742.PLACE_LOCATION = "NONE";
      defparam ii3742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3743 ( .DX(nn3743), .F0(nn3655), .F1(dummy_431_), .F2(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ), .F3(dummy_abc_2590_) );
      defparam ii3743.CONFIG_DATA = 16'hB8B8;
      defparam ii3743.PLACE_LOCATION = "NONE";
      defparam ii3743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3744 ( .DX(nn3744), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2591_), .F3(dummy_abc_2592_) );
      defparam ii3744.CONFIG_DATA = 16'h9999;
      defparam ii3744.PLACE_LOCATION = "NONE";
      defparam ii3744.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3745 ( .DX(nn3745), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_431_) );
      defparam ii3745.CONFIG_DATA = 16'hA569;
      defparam ii3745.PLACE_LOCATION = "NONE";
      defparam ii3745.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3746 ( .DX(nn3746), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_431_), .F2(nn3645), .F3(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ) );
      defparam ii3746.CONFIG_DATA = 16'hA695;
      defparam ii3746.PLACE_LOCATION = "NONE";
      defparam ii3746.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3747 ( .DX(nn3747), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3646), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ) );
      defparam ii3747.CONFIG_DATA = 16'h9A95;
      defparam ii3747.PLACE_LOCATION = "NONE";
      defparam ii3747.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3748 ( .DX(nn3748), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3647), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ) );
      defparam ii3748.CONFIG_DATA = 16'h9A95;
      defparam ii3748.PLACE_LOCATION = "NONE";
      defparam ii3748.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3749 ( .DX(nn3749), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3648), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ) );
      defparam ii3749.CONFIG_DATA = 16'h9A95;
      defparam ii3749.PLACE_LOCATION = "NONE";
      defparam ii3749.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3750 ( .DX(nn3750), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3649), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ) );
      defparam ii3750.CONFIG_DATA = 16'h9A95;
      defparam ii3750.PLACE_LOCATION = "NONE";
      defparam ii3750.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3751 ( .DX(nn3751), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3650), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ) );
      defparam ii3751.CONFIG_DATA = 16'h9A95;
      defparam ii3751.PLACE_LOCATION = "NONE";
      defparam ii3751.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3752 ( .DX(nn3752), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3651), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ) );
      defparam ii3752.CONFIG_DATA = 16'h9A95;
      defparam ii3752.PLACE_LOCATION = "NONE";
      defparam ii3752.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3753 ( .DX(nn3753), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3652), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ) );
      defparam ii3753.CONFIG_DATA = 16'h9A95;
      defparam ii3753.PLACE_LOCATION = "NONE";
      defparam ii3753.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3754 ( .DX(nn3754), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3653), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ) );
      defparam ii3754.CONFIG_DATA = 16'h9A95;
      defparam ii3754.PLACE_LOCATION = "NONE";
      defparam ii3754.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3755 ( .DX(nn3755), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3654), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ) );
      defparam ii3755.CONFIG_DATA = 16'h9A95;
      defparam ii3755.PLACE_LOCATION = "NONE";
      defparam ii3755.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3756 ( .DX(nn3756), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3655), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ) );
      defparam ii3756.CONFIG_DATA = 16'h9A95;
      defparam ii3756.PLACE_LOCATION = "NONE";
      defparam ii3756.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3757 ( .DX(nn3757), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3706), .F2(dummy_431_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3757.CONFIG_DATA = 16'h9095;
      defparam ii3757.PLACE_LOCATION = "NONE";
      defparam ii3757.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3758 ( .DX(nn3758), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2593_), .F2(dummy_abc_2594_), .F3(dummy_abc_2595_) );
      defparam ii3758.CONFIG_DATA = 16'h5555;
      defparam ii3758.PLACE_LOCATION = "NONE";
      defparam ii3758.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3759 ( .DX(nn3759), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2596_), .F2(dummy_abc_2597_), .F3(dummy_abc_2598_) );
      defparam ii3759.CONFIG_DATA = 16'h5555;
      defparam ii3759.PLACE_LOCATION = "NONE";
      defparam ii3759.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3760 ( .DX(nn3760), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2599_), .F2(dummy_abc_2600_), .F3(dummy_abc_2601_) );
      defparam ii3760.CONFIG_DATA = 16'h5555;
      defparam ii3760.PLACE_LOCATION = "NONE";
      defparam ii3760.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_21_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, nn3692, nn3743, nn3742, nn3741, nn3740, nn3739, nn3738, 
              nn3737, nn3736, nn3735, nn3734, nn3733, nn3732, 
              \coefcal1_xDividend__reg[3]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_162_ ), 
        .DX( {nn3760, nn3759, nn3758, nn3757, nn3756, nn3755, nn3754, nn3753, 
              nn3752, nn3751, nn3750, nn3749, nn3748, nn3747, nn3746, nn3745, 
              nn3744} ), 
        .SUM( {dummy_163_, \coefcal1_divide_inst1_u114_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_14|SUM_net , \coefcal1_divide_inst1_u114_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_12|SUM_net , \coefcal1_divide_inst1_u114_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_10|SUM_net , \coefcal1_divide_inst1_u114_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_8|SUM_net , \coefcal1_divide_inst1_u114_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_6|SUM_net , \coefcal1_divide_inst1_u114_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_4|SUM_net , \coefcal1_divide_inst1_u114_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_2|SUM_net , \coefcal1_divide_inst1_u114_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3780 ( .DX(nn3780), .F0(nn3692), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ), .F3(dummy_abc_2602_) );
      defparam ii3780.CONFIG_DATA = 16'hA8A8;
      defparam ii3780.PLACE_LOCATION = "NONE";
      defparam ii3780.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3781 ( .DX(nn3781), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2603_), .F3(dummy_abc_2604_) );
      defparam ii3781.CONFIG_DATA = 16'h9999;
      defparam ii3781.PLACE_LOCATION = "NONE";
      defparam ii3781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3782 ( .DX(nn3782), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_450_) );
      defparam ii3782.CONFIG_DATA = 16'hA569;
      defparam ii3782.PLACE_LOCATION = "NONE";
      defparam ii3782.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3783 ( .DX(nn3783), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_450_), .F2(nn3732), .F3(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ) );
      defparam ii3783.CONFIG_DATA = 16'hA695;
      defparam ii3783.PLACE_LOCATION = "NONE";
      defparam ii3783.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3784 ( .DX(nn3784), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3733), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ) );
      defparam ii3784.CONFIG_DATA = 16'h9A95;
      defparam ii3784.PLACE_LOCATION = "NONE";
      defparam ii3784.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3785 ( .DX(nn3785), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3734), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ) );
      defparam ii3785.CONFIG_DATA = 16'h9A95;
      defparam ii3785.PLACE_LOCATION = "NONE";
      defparam ii3785.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3786 ( .DX(nn3786), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3735), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ) );
      defparam ii3786.CONFIG_DATA = 16'h9A95;
      defparam ii3786.PLACE_LOCATION = "NONE";
      defparam ii3786.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3787 ( .DX(nn3787), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3736), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ) );
      defparam ii3787.CONFIG_DATA = 16'h9A95;
      defparam ii3787.PLACE_LOCATION = "NONE";
      defparam ii3787.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3788 ( .DX(nn3788), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3737), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ) );
      defparam ii3788.CONFIG_DATA = 16'h9A95;
      defparam ii3788.PLACE_LOCATION = "NONE";
      defparam ii3788.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3789 ( .DX(nn3789), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3738), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ) );
      defparam ii3789.CONFIG_DATA = 16'h9A95;
      defparam ii3789.PLACE_LOCATION = "NONE";
      defparam ii3789.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3790 ( .DX(nn3790), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3739), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ) );
      defparam ii3790.CONFIG_DATA = 16'h9A95;
      defparam ii3790.PLACE_LOCATION = "NONE";
      defparam ii3790.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3791 ( .DX(nn3791), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3740), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ) );
      defparam ii3791.CONFIG_DATA = 16'h9A95;
      defparam ii3791.PLACE_LOCATION = "NONE";
      defparam ii3791.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3792 ( .DX(nn3792), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3741), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ) );
      defparam ii3792.CONFIG_DATA = 16'h9A95;
      defparam ii3792.PLACE_LOCATION = "NONE";
      defparam ii3792.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3793 ( .DX(nn3793), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3742), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ) );
      defparam ii3793.CONFIG_DATA = 16'h9A95;
      defparam ii3793.PLACE_LOCATION = "NONE";
      defparam ii3793.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3794 ( .DX(nn3794), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3743), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ) );
      defparam ii3794.CONFIG_DATA = 16'h9A95;
      defparam ii3794.PLACE_LOCATION = "NONE";
      defparam ii3794.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3795 ( .DX(nn3795), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3692), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ) );
      defparam ii3795.CONFIG_DATA = 16'h9995;
      defparam ii3795.PLACE_LOCATION = "NONE";
      defparam ii3795.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3796 ( .DX(nn3796), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2605_), .F2(dummy_abc_2606_), .F3(dummy_abc_2607_) );
      defparam ii3796.CONFIG_DATA = 16'h5555;
      defparam ii3796.PLACE_LOCATION = "NONE";
      defparam ii3796.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3797 ( .DX(nn3797), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2608_), .F2(dummy_abc_2609_), .F3(dummy_abc_2610_) );
      defparam ii3797.CONFIG_DATA = 16'h5555;
      defparam ii3797.PLACE_LOCATION = "NONE";
      defparam ii3797.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3798 ( .DX(nn3798), .F0(dummy_abc_2611_), .F1(dummy_abc_2612_), .F2(dummy_abc_2613_), .F3(dummy_abc_2614_) );
      defparam ii3798.CONFIG_DATA = 16'hFFFF;
      defparam ii3798.PLACE_LOCATION = "NONE";
      defparam ii3798.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_37_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_469_ ), 
        .DX( {nn3798, nn3797, nn3796, nn3795, nn3794, nn3793, nn3792, nn3791, 
              nn3790, nn3789, nn3788, nn3787, nn3786, nn3785, nn3784, nn3783, 
              nn3782, nn3781} ), 
        .SUM( {\coefcal1_divide_inst1_u146_XORCI_17|SUM_net , dummy_470_, 
              dummy_471_, dummy_472_, dummy_473_, dummy_474_, dummy_475_, dummy_476_, 
              dummy_477_, dummy_478_, dummy_479_, dummy_480_, dummy_481_, dummy_482_, 
              dummy_483_, dummy_484_, dummy_485_, dummy_486_} )
      );
    CS_LUT4_PRIM ii3819 ( .DX(nn3819), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_450_), .F3(dummy_abc_2615_) );
      defparam ii3819.CONFIG_DATA = 16'hA6A6;
      defparam ii3819.PLACE_LOCATION = "NONE";
      defparam ii3819.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3820 ( .DX(nn3820), .F0(dummy_450_), .F1(nn3732), .F2(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ), .F3(dummy_abc_2616_) );
      defparam ii3820.CONFIG_DATA = 16'hD8D8;
      defparam ii3820.PLACE_LOCATION = "NONE";
      defparam ii3820.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3821 ( .DX(nn3821), .F0(nn3733), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ), .F3(dummy_abc_2617_) );
      defparam ii3821.CONFIG_DATA = 16'hB8B8;
      defparam ii3821.PLACE_LOCATION = "NONE";
      defparam ii3821.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3822 ( .DX(nn3822), .F0(nn3734), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ), .F3(dummy_abc_2618_) );
      defparam ii3822.CONFIG_DATA = 16'hB8B8;
      defparam ii3822.PLACE_LOCATION = "NONE";
      defparam ii3822.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3823 ( .DX(nn3823), .F0(nn3735), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ), .F3(dummy_abc_2619_) );
      defparam ii3823.CONFIG_DATA = 16'hB8B8;
      defparam ii3823.PLACE_LOCATION = "NONE";
      defparam ii3823.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3824 ( .DX(nn3824), .F0(nn3736), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ), .F3(dummy_abc_2620_) );
      defparam ii3824.CONFIG_DATA = 16'hB8B8;
      defparam ii3824.PLACE_LOCATION = "NONE";
      defparam ii3824.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3825 ( .DX(nn3825), .F0(nn3737), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ), .F3(dummy_abc_2621_) );
      defparam ii3825.CONFIG_DATA = 16'hB8B8;
      defparam ii3825.PLACE_LOCATION = "NONE";
      defparam ii3825.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3826 ( .DX(nn3826), .F0(nn3738), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ), .F3(dummy_abc_2622_) );
      defparam ii3826.CONFIG_DATA = 16'hB8B8;
      defparam ii3826.PLACE_LOCATION = "NONE";
      defparam ii3826.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3827 ( .DX(nn3827), .F0(nn3739), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ), .F3(dummy_abc_2623_) );
      defparam ii3827.CONFIG_DATA = 16'hB8B8;
      defparam ii3827.PLACE_LOCATION = "NONE";
      defparam ii3827.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3828 ( .DX(nn3828), .F0(nn3740), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ), .F3(dummy_abc_2624_) );
      defparam ii3828.CONFIG_DATA = 16'hB8B8;
      defparam ii3828.PLACE_LOCATION = "NONE";
      defparam ii3828.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3829 ( .DX(nn3829), .F0(nn3741), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ), .F3(dummy_abc_2625_) );
      defparam ii3829.CONFIG_DATA = 16'hB8B8;
      defparam ii3829.PLACE_LOCATION = "NONE";
      defparam ii3829.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3830 ( .DX(nn3830), .F0(nn3742), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ), .F3(dummy_abc_2626_) );
      defparam ii3830.CONFIG_DATA = 16'hB8B8;
      defparam ii3830.PLACE_LOCATION = "NONE";
      defparam ii3830.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3831 ( .DX(nn3831), .F0(nn3743), .F1(dummy_450_), .F2(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ), .F3(dummy_abc_2627_) );
      defparam ii3831.CONFIG_DATA = 16'hB8B8;
      defparam ii3831.PLACE_LOCATION = "NONE";
      defparam ii3831.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3832 ( .DX(nn3832), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2628_), .F3(dummy_abc_2629_) );
      defparam ii3832.CONFIG_DATA = 16'h9999;
      defparam ii3832.PLACE_LOCATION = "NONE";
      defparam ii3832.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3833 ( .DX(nn3833), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_450_) );
      defparam ii3833.CONFIG_DATA = 16'hA569;
      defparam ii3833.PLACE_LOCATION = "NONE";
      defparam ii3833.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3834 ( .DX(nn3834), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_450_), .F2(nn3732), .F3(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ) );
      defparam ii3834.CONFIG_DATA = 16'hA695;
      defparam ii3834.PLACE_LOCATION = "NONE";
      defparam ii3834.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3835 ( .DX(nn3835), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3733), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ) );
      defparam ii3835.CONFIG_DATA = 16'h9A95;
      defparam ii3835.PLACE_LOCATION = "NONE";
      defparam ii3835.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3836 ( .DX(nn3836), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3734), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ) );
      defparam ii3836.CONFIG_DATA = 16'h9A95;
      defparam ii3836.PLACE_LOCATION = "NONE";
      defparam ii3836.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3837 ( .DX(nn3837), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3735), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ) );
      defparam ii3837.CONFIG_DATA = 16'h9A95;
      defparam ii3837.PLACE_LOCATION = "NONE";
      defparam ii3837.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3838 ( .DX(nn3838), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3736), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ) );
      defparam ii3838.CONFIG_DATA = 16'h9A95;
      defparam ii3838.PLACE_LOCATION = "NONE";
      defparam ii3838.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3839 ( .DX(nn3839), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3737), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ) );
      defparam ii3839.CONFIG_DATA = 16'h9A95;
      defparam ii3839.PLACE_LOCATION = "NONE";
      defparam ii3839.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3840 ( .DX(nn3840), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3738), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ) );
      defparam ii3840.CONFIG_DATA = 16'h9A95;
      defparam ii3840.PLACE_LOCATION = "NONE";
      defparam ii3840.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3841 ( .DX(nn3841), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3739), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ) );
      defparam ii3841.CONFIG_DATA = 16'h9A95;
      defparam ii3841.PLACE_LOCATION = "NONE";
      defparam ii3841.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3842 ( .DX(nn3842), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3740), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ) );
      defparam ii3842.CONFIG_DATA = 16'h9A95;
      defparam ii3842.PLACE_LOCATION = "NONE";
      defparam ii3842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3843 ( .DX(nn3843), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3741), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ) );
      defparam ii3843.CONFIG_DATA = 16'h9A95;
      defparam ii3843.PLACE_LOCATION = "NONE";
      defparam ii3843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3844 ( .DX(nn3844), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3742), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ) );
      defparam ii3844.CONFIG_DATA = 16'h9A95;
      defparam ii3844.PLACE_LOCATION = "NONE";
      defparam ii3844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3845 ( .DX(nn3845), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3743), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ) );
      defparam ii3845.CONFIG_DATA = 16'h9A95;
      defparam ii3845.PLACE_LOCATION = "NONE";
      defparam ii3845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3846 ( .DX(nn3846), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3692), .F2(dummy_450_), .F3(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ) );
      defparam ii3846.CONFIG_DATA = 16'h9995;
      defparam ii3846.PLACE_LOCATION = "NONE";
      defparam ii3846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3847 ( .DX(nn3847), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2630_), .F2(dummy_abc_2631_), .F3(dummy_abc_2632_) );
      defparam ii3847.CONFIG_DATA = 16'h5555;
      defparam ii3847.PLACE_LOCATION = "NONE";
      defparam ii3847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3848 ( .DX(nn3848), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2633_), .F2(dummy_abc_2634_), .F3(dummy_abc_2635_) );
      defparam ii3848.CONFIG_DATA = 16'h5555;
      defparam ii3848.PLACE_LOCATION = "NONE";
      defparam ii3848.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_22_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, nn3780, nn3831, 
              nn3830, nn3829, nn3828, nn3827, nn3826, nn3825, nn3824, nn3823, 
              nn3822, nn3821, nn3820, nn3819, \coefcal1_xDividend__reg[2]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_164_ ), 
        .DX( {nn3848, nn3847, nn3846, nn3845, nn3844, nn3843, nn3842, nn3841, 
              nn3840, nn3839, nn3838, nn3837, nn3836, nn3835, nn3834, nn3833, 
              nn3832} ), 
        .SUM( {dummy_165_, \coefcal1_divide_inst1_u115_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_14|SUM_net , \coefcal1_divide_inst1_u115_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_12|SUM_net , \coefcal1_divide_inst1_u115_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_10|SUM_net , \coefcal1_divide_inst1_u115_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_8|SUM_net , \coefcal1_divide_inst1_u115_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_6|SUM_net , \coefcal1_divide_inst1_u115_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_4|SUM_net , \coefcal1_divide_inst1_u115_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_2|SUM_net , \coefcal1_divide_inst1_u115_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3868 ( .DX(nn3868), .F0(nn3780), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_14|SUM_net ), .F3(dummy_abc_2636_) );
      defparam ii3868.CONFIG_DATA = 16'hB8B8;
      defparam ii3868.PLACE_LOCATION = "NONE";
      defparam ii3868.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3869 ( .DX(nn3869), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2637_), .F3(dummy_abc_2638_) );
      defparam ii3869.CONFIG_DATA = 16'h9999;
      defparam ii3869.PLACE_LOCATION = "NONE";
      defparam ii3869.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3870 ( .DX(nn3870), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_469_) );
      defparam ii3870.CONFIG_DATA = 16'hA569;
      defparam ii3870.PLACE_LOCATION = "NONE";
      defparam ii3870.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3871 ( .DX(nn3871), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_469_), .F2(nn3819), .F3(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ) );
      defparam ii3871.CONFIG_DATA = 16'hA695;
      defparam ii3871.PLACE_LOCATION = "NONE";
      defparam ii3871.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3872 ( .DX(nn3872), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3820), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_2|SUM_net ) );
      defparam ii3872.CONFIG_DATA = 16'h9A95;
      defparam ii3872.PLACE_LOCATION = "NONE";
      defparam ii3872.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3873 ( .DX(nn3873), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3821), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_3|SUM_net ) );
      defparam ii3873.CONFIG_DATA = 16'h9A95;
      defparam ii3873.PLACE_LOCATION = "NONE";
      defparam ii3873.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3874 ( .DX(nn3874), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3822), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_4|SUM_net ) );
      defparam ii3874.CONFIG_DATA = 16'h9A95;
      defparam ii3874.PLACE_LOCATION = "NONE";
      defparam ii3874.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3875 ( .DX(nn3875), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3823), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_5|SUM_net ) );
      defparam ii3875.CONFIG_DATA = 16'h9A95;
      defparam ii3875.PLACE_LOCATION = "NONE";
      defparam ii3875.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3876 ( .DX(nn3876), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3824), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_6|SUM_net ) );
      defparam ii3876.CONFIG_DATA = 16'h9A95;
      defparam ii3876.PLACE_LOCATION = "NONE";
      defparam ii3876.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3877 ( .DX(nn3877), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3825), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_7|SUM_net ) );
      defparam ii3877.CONFIG_DATA = 16'h9A95;
      defparam ii3877.PLACE_LOCATION = "NONE";
      defparam ii3877.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3878 ( .DX(nn3878), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3826), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_8|SUM_net ) );
      defparam ii3878.CONFIG_DATA = 16'h9A95;
      defparam ii3878.PLACE_LOCATION = "NONE";
      defparam ii3878.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3879 ( .DX(nn3879), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3827), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_9|SUM_net ) );
      defparam ii3879.CONFIG_DATA = 16'h9A95;
      defparam ii3879.PLACE_LOCATION = "NONE";
      defparam ii3879.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3880 ( .DX(nn3880), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3828), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_10|SUM_net ) );
      defparam ii3880.CONFIG_DATA = 16'h9A95;
      defparam ii3880.PLACE_LOCATION = "NONE";
      defparam ii3880.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3881 ( .DX(nn3881), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3829), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_11|SUM_net ) );
      defparam ii3881.CONFIG_DATA = 16'h9A95;
      defparam ii3881.PLACE_LOCATION = "NONE";
      defparam ii3881.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3882 ( .DX(nn3882), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3830), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_12|SUM_net ) );
      defparam ii3882.CONFIG_DATA = 16'h9A95;
      defparam ii3882.PLACE_LOCATION = "NONE";
      defparam ii3882.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3883 ( .DX(nn3883), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3831), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_13|SUM_net ) );
      defparam ii3883.CONFIG_DATA = 16'h9A95;
      defparam ii3883.PLACE_LOCATION = "NONE";
      defparam ii3883.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3884 ( .DX(nn3884), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn3780), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_14|SUM_net ) );
      defparam ii3884.CONFIG_DATA = 16'h9A95;
      defparam ii3884.PLACE_LOCATION = "NONE";
      defparam ii3884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3885 ( .DX(nn3885), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2639_), .F2(dummy_abc_2640_), .F3(dummy_abc_2641_) );
      defparam ii3885.CONFIG_DATA = 16'h5555;
      defparam ii3885.PLACE_LOCATION = "NONE";
      defparam ii3885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3886 ( .DX(nn3886), .F0(dummy_abc_2642_), .F1(dummy_abc_2643_), .F2(dummy_abc_2644_), .F3(dummy_abc_2645_) );
      defparam ii3886.CONFIG_DATA = 16'hFFFF;
      defparam ii3886.PLACE_LOCATION = "NONE";
      defparam ii3886.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_38_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_488_ ), 
        .DX( {nn3886, nn3885, nn3884, nn3883, nn3882, nn3881, nn3880, nn3879, 
              nn3878, nn3877, nn3876, nn3875, nn3874, nn3873, nn3872, nn3871, 
              nn3870, nn3869} ), 
        .SUM( {\coefcal1_divide_inst1_u148_XORCI_17|SUM_net , dummy_489_, 
              dummy_490_, dummy_491_, dummy_492_, dummy_493_, dummy_494_, dummy_495_, 
              dummy_496_, dummy_497_, dummy_498_, dummy_499_, dummy_500_, dummy_501_, 
              dummy_502_, dummy_503_, dummy_504_, dummy_505_} )
      );
    CS_LUT4_PRIM ii3907 ( .DX(nn3907), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_469_), .F3(dummy_abc_2646_) );
      defparam ii3907.CONFIG_DATA = 16'hA6A6;
      defparam ii3907.PLACE_LOCATION = "NONE";
      defparam ii3907.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3908 ( .DX(nn3908), .F0(dummy_469_), .F1(nn3819), .F2(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ), .F3(dummy_abc_2647_) );
      defparam ii3908.CONFIG_DATA = 16'hD8D8;
      defparam ii3908.PLACE_LOCATION = "NONE";
      defparam ii3908.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3909 ( .DX(nn3909), .F0(nn3820), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_2|SUM_net ), .F3(dummy_abc_2648_) );
      defparam ii3909.CONFIG_DATA = 16'hB8B8;
      defparam ii3909.PLACE_LOCATION = "NONE";
      defparam ii3909.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3910 ( .DX(nn3910), .F0(nn3821), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_3|SUM_net ), .F3(dummy_abc_2649_) );
      defparam ii3910.CONFIG_DATA = 16'hB8B8;
      defparam ii3910.PLACE_LOCATION = "NONE";
      defparam ii3910.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3911 ( .DX(nn3911), .F0(nn3822), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_4|SUM_net ), .F3(dummy_abc_2650_) );
      defparam ii3911.CONFIG_DATA = 16'hB8B8;
      defparam ii3911.PLACE_LOCATION = "NONE";
      defparam ii3911.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3912 ( .DX(nn3912), .F0(nn3823), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_5|SUM_net ), .F3(dummy_abc_2651_) );
      defparam ii3912.CONFIG_DATA = 16'hB8B8;
      defparam ii3912.PLACE_LOCATION = "NONE";
      defparam ii3912.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3913 ( .DX(nn3913), .F0(nn3824), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_6|SUM_net ), .F3(dummy_abc_2652_) );
      defparam ii3913.CONFIG_DATA = 16'hB8B8;
      defparam ii3913.PLACE_LOCATION = "NONE";
      defparam ii3913.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3914 ( .DX(nn3914), .F0(nn3825), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_7|SUM_net ), .F3(dummy_abc_2653_) );
      defparam ii3914.CONFIG_DATA = 16'hB8B8;
      defparam ii3914.PLACE_LOCATION = "NONE";
      defparam ii3914.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3915 ( .DX(nn3915), .F0(nn3826), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_8|SUM_net ), .F3(dummy_abc_2654_) );
      defparam ii3915.CONFIG_DATA = 16'hB8B8;
      defparam ii3915.PLACE_LOCATION = "NONE";
      defparam ii3915.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3916 ( .DX(nn3916), .F0(nn3827), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_9|SUM_net ), .F3(dummy_abc_2655_) );
      defparam ii3916.CONFIG_DATA = 16'hB8B8;
      defparam ii3916.PLACE_LOCATION = "NONE";
      defparam ii3916.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3917 ( .DX(nn3917), .F0(nn3828), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_10|SUM_net ), .F3(dummy_abc_2656_) );
      defparam ii3917.CONFIG_DATA = 16'hB8B8;
      defparam ii3917.PLACE_LOCATION = "NONE";
      defparam ii3917.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3918 ( .DX(nn3918), .F0(nn3829), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_11|SUM_net ), .F3(dummy_abc_2657_) );
      defparam ii3918.CONFIG_DATA = 16'hB8B8;
      defparam ii3918.PLACE_LOCATION = "NONE";
      defparam ii3918.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3919 ( .DX(nn3919), .F0(nn3830), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_12|SUM_net ), .F3(dummy_abc_2658_) );
      defparam ii3919.CONFIG_DATA = 16'hB8B8;
      defparam ii3919.PLACE_LOCATION = "NONE";
      defparam ii3919.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3920 ( .DX(nn3920), .F0(nn3831), .F1(dummy_469_), .F2(\coefcal1_divide_inst1_u115_XORCI_13|SUM_net ), .F3(dummy_abc_2659_) );
      defparam ii3920.CONFIG_DATA = 16'hB8B8;
      defparam ii3920.PLACE_LOCATION = "NONE";
      defparam ii3920.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3921 ( .DX(nn3921), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2660_), .F3(dummy_abc_2661_) );
      defparam ii3921.CONFIG_DATA = 16'h9999;
      defparam ii3921.PLACE_LOCATION = "NONE";
      defparam ii3921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3922 ( .DX(nn3922), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_469_) );
      defparam ii3922.CONFIG_DATA = 16'hA569;
      defparam ii3922.PLACE_LOCATION = "NONE";
      defparam ii3922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3923 ( .DX(nn3923), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_469_), .F2(nn3819), .F3(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ) );
      defparam ii3923.CONFIG_DATA = 16'hA695;
      defparam ii3923.PLACE_LOCATION = "NONE";
      defparam ii3923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3924 ( .DX(nn3924), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3820), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_2|SUM_net ) );
      defparam ii3924.CONFIG_DATA = 16'h9A95;
      defparam ii3924.PLACE_LOCATION = "NONE";
      defparam ii3924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3925 ( .DX(nn3925), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3821), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_3|SUM_net ) );
      defparam ii3925.CONFIG_DATA = 16'h9A95;
      defparam ii3925.PLACE_LOCATION = "NONE";
      defparam ii3925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3926 ( .DX(nn3926), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3822), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_4|SUM_net ) );
      defparam ii3926.CONFIG_DATA = 16'h9A95;
      defparam ii3926.PLACE_LOCATION = "NONE";
      defparam ii3926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3927 ( .DX(nn3927), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3823), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_5|SUM_net ) );
      defparam ii3927.CONFIG_DATA = 16'h9A95;
      defparam ii3927.PLACE_LOCATION = "NONE";
      defparam ii3927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3928 ( .DX(nn3928), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3824), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_6|SUM_net ) );
      defparam ii3928.CONFIG_DATA = 16'h9A95;
      defparam ii3928.PLACE_LOCATION = "NONE";
      defparam ii3928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3929 ( .DX(nn3929), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3825), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_7|SUM_net ) );
      defparam ii3929.CONFIG_DATA = 16'h9A95;
      defparam ii3929.PLACE_LOCATION = "NONE";
      defparam ii3929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3930 ( .DX(nn3930), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3826), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_8|SUM_net ) );
      defparam ii3930.CONFIG_DATA = 16'h9A95;
      defparam ii3930.PLACE_LOCATION = "NONE";
      defparam ii3930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3931 ( .DX(nn3931), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3827), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_9|SUM_net ) );
      defparam ii3931.CONFIG_DATA = 16'h9A95;
      defparam ii3931.PLACE_LOCATION = "NONE";
      defparam ii3931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3932 ( .DX(nn3932), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3828), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_10|SUM_net ) );
      defparam ii3932.CONFIG_DATA = 16'h9A95;
      defparam ii3932.PLACE_LOCATION = "NONE";
      defparam ii3932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3933 ( .DX(nn3933), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3829), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_11|SUM_net ) );
      defparam ii3933.CONFIG_DATA = 16'h9A95;
      defparam ii3933.PLACE_LOCATION = "NONE";
      defparam ii3933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3934 ( .DX(nn3934), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3830), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_12|SUM_net ) );
      defparam ii3934.CONFIG_DATA = 16'h9A95;
      defparam ii3934.PLACE_LOCATION = "NONE";
      defparam ii3934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3935 ( .DX(nn3935), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3831), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_13|SUM_net ) );
      defparam ii3935.CONFIG_DATA = 16'h9A95;
      defparam ii3935.PLACE_LOCATION = "NONE";
      defparam ii3935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3936 ( .DX(nn3936), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn3780), .F2(dummy_469_), .F3(\coefcal1_divide_inst1_u115_XORCI_14|SUM_net ) );
      defparam ii3936.CONFIG_DATA = 16'h9A95;
      defparam ii3936.PLACE_LOCATION = "NONE";
      defparam ii3936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3937 ( .DX(nn3937), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2662_), .F2(dummy_abc_2663_), .F3(dummy_abc_2664_) );
      defparam ii3937.CONFIG_DATA = 16'h5555;
      defparam ii3937.PLACE_LOCATION = "NONE";
      defparam ii3937.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_23_ ( 
        .CA( {a_acc_en_cal1_u134_mac, nn3868, nn3920, nn3919, nn3918, nn3917, 
              nn3916, nn3915, nn3914, nn3913, nn3912, nn3911, nn3910, nn3909, 
              nn3908, nn3907, \coefcal1_xDividend__reg[1]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_166_ ), 
        .DX( {nn3937, nn3936, nn3935, nn3934, nn3933, nn3932, nn3931, nn3930, 
              nn3929, nn3928, nn3927, nn3926, nn3925, nn3924, nn3923, nn3922, 
              nn3921} ), 
        .SUM( {dummy_167_, \coefcal1_divide_inst1_u116_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_14|SUM_net , \coefcal1_divide_inst1_u116_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_12|SUM_net , \coefcal1_divide_inst1_u116_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_10|SUM_net , \coefcal1_divide_inst1_u116_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_8|SUM_net , \coefcal1_divide_inst1_u116_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_6|SUM_net , \coefcal1_divide_inst1_u116_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_4|SUM_net , \coefcal1_divide_inst1_u116_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_2|SUM_net , \coefcal1_divide_inst1_u116_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3957 ( .DX(nn3957), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(nn3868), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_15|SUM_net ) );
      defparam ii3957.CONFIG_DATA = 16'h8A80;
      defparam ii3957.PLACE_LOCATION = "NONE";
      defparam ii3957.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3958 ( .DX(nn3958), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[16]|Q_net ), .F2(nn3957), .F3(dummy_abc_2665_) );
      defparam ii3958.CONFIG_DATA = 16'hF1F1;
      defparam ii3958.PLACE_LOCATION = "NONE";
      defparam ii3958.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3959 ( .DX(nn3959), .F0(dummy_abc_2666_), .F1(dummy_abc_2667_), .F2(dummy_abc_2668_), .F3(dummy_abc_2669_) );
      defparam ii3959.CONFIG_DATA = 16'hFFFF;
      defparam ii3959.PLACE_LOCATION = "NONE";
      defparam ii3959.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18 ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDividend__reg[16]|Q_net , 
              \coefcal1_xDividend__reg[15]|Q_net , \coefcal1_xDividend__reg[14]|Q_net , 
              \coefcal1_xDividend__reg[13]|Q_net , \coefcal1_xDividend__reg[12]|Q_net , 
              \coefcal1_xDividend__reg[11]|Q_net , \coefcal1_xDividend__reg[10]|Q_net , 
              \coefcal1_xDividend__reg[9]|Q_net , \coefcal1_xDividend__reg[8]|Q_net , 
              \coefcal1_xDividend__reg[7]|Q_net , \coefcal1_xDividend__reg[6]|Q_net , 
              \coefcal1_xDividend__reg[5]|Q_net , \coefcal1_xDividend__reg[4]|Q_net , 
              \coefcal1_xDividend__reg[3]|Q_net , \coefcal1_xDividend__reg[2]|Q_net , 
              \coefcal1_xDividend__reg[1]|Q_net , \coefcal1_xDividend__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_203_ ), 
        .DX( {nn3959, nn3958, nn2727, nn2726, nn2725, nn2724, nn2723, nn2722, 
              nn2721, nn2720, nn2719, nn2718, nn2717, nn2716, nn2715, nn2714, 
              nn2713, nn2712} ), 
        .SUM( {\coefcal1_divide_inst1_u118_XORCI_17|SUM_net , dummy_204_, 
              dummy_205_, dummy_206_, dummy_207_, dummy_208_, dummy_209_, dummy_210_, 
              dummy_211_, dummy_212_, dummy_213_, dummy_214_, dummy_215_, dummy_216_, 
              dummy_217_, dummy_218_, dummy_219_, dummy_220_} )
      );
    CS_LUT4_PRIM ii3980 ( .DX(nn3980), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[15]|Q_net ), .F2(\coefcal1_xDivisor__reg[16]|Q_net ), .F3(\coefcal1_xDivisor__reg[1]|Q_net ) );
      defparam ii3980.CONFIG_DATA = 16'h0001;
      defparam ii3980.PLACE_LOCATION = "NONE";
      defparam ii3980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3981 ( .DX(nn3981), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[11]|Q_net ), .F2(\coefcal1_xDivisor__reg[12]|Q_net ), .F3(nn3980) );
      defparam ii3981.CONFIG_DATA = 16'h0100;
      defparam ii3981.PLACE_LOCATION = "NONE";
      defparam ii3981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3982 ( .DX(nn3982), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[7]|Q_net ), .F2(\coefcal1_xDivisor__reg[8]|Q_net ), .F3(\coefcal1_xDivisor__reg[9]|Q_net ) );
      defparam ii3982.CONFIG_DATA = 16'h0001;
      defparam ii3982.PLACE_LOCATION = "NONE";
      defparam ii3982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3983 ( .DX(nn3983), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[3]|Q_net ), .F2(\coefcal1_xDivisor__reg[5]|Q_net ), .F3(nn3982) );
      defparam ii3983.CONFIG_DATA = 16'h0100;
      defparam ii3983.PLACE_LOCATION = "NONE";
      defparam ii3983.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3984 ( .DX(nn3984), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[4]|Q_net ), .F2(nn3981), .F3(nn3983) );
      defparam ii3984.CONFIG_DATA = 16'h1000;
      defparam ii3984.PLACE_LOCATION = "NONE";
      defparam ii3984.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3985 ( .DX(nn3985), .F0(\coefcal1_xDivisor__reg[0]|Q_net ), .F1(nn3984), .F2(dummy_abc_2670_), .F3(dummy_abc_2671_) );
      defparam ii3985.CONFIG_DATA = 16'h4444;
      defparam ii3985.PLACE_LOCATION = "NONE";
      defparam ii3985.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3986 ( .DX(nn3986), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2672_), .F3(dummy_abc_2673_) );
      defparam ii3986.CONFIG_DATA = 16'h9999;
      defparam ii3986.PLACE_LOCATION = "NONE";
      defparam ii3986.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3987 ( .DX(nn3987), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_488_) );
      defparam ii3987.CONFIG_DATA = 16'hA569;
      defparam ii3987.PLACE_LOCATION = "NONE";
      defparam ii3987.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3988 ( .DX(nn3988), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_488_), .F2(nn3907), .F3(\coefcal1_divide_inst1_u116_XORCI_1|SUM_net ) );
      defparam ii3988.CONFIG_DATA = 16'hA695;
      defparam ii3988.PLACE_LOCATION = "NONE";
      defparam ii3988.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3989 ( .DX(nn3989), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3908), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_2|SUM_net ) );
      defparam ii3989.CONFIG_DATA = 16'h9A95;
      defparam ii3989.PLACE_LOCATION = "NONE";
      defparam ii3989.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3990 ( .DX(nn3990), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3909), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_3|SUM_net ) );
      defparam ii3990.CONFIG_DATA = 16'h9A95;
      defparam ii3990.PLACE_LOCATION = "NONE";
      defparam ii3990.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3991 ( .DX(nn3991), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3910), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_4|SUM_net ) );
      defparam ii3991.CONFIG_DATA = 16'h9A95;
      defparam ii3991.PLACE_LOCATION = "NONE";
      defparam ii3991.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3992 ( .DX(nn3992), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3911), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_5|SUM_net ) );
      defparam ii3992.CONFIG_DATA = 16'h9A95;
      defparam ii3992.PLACE_LOCATION = "NONE";
      defparam ii3992.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3993 ( .DX(nn3993), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3912), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_6|SUM_net ) );
      defparam ii3993.CONFIG_DATA = 16'h9A95;
      defparam ii3993.PLACE_LOCATION = "NONE";
      defparam ii3993.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3994 ( .DX(nn3994), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3913), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_7|SUM_net ) );
      defparam ii3994.CONFIG_DATA = 16'h9A95;
      defparam ii3994.PLACE_LOCATION = "NONE";
      defparam ii3994.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3995 ( .DX(nn3995), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3914), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_8|SUM_net ) );
      defparam ii3995.CONFIG_DATA = 16'h9A95;
      defparam ii3995.PLACE_LOCATION = "NONE";
      defparam ii3995.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3996 ( .DX(nn3996), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3915), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_9|SUM_net ) );
      defparam ii3996.CONFIG_DATA = 16'h9A95;
      defparam ii3996.PLACE_LOCATION = "NONE";
      defparam ii3996.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3997 ( .DX(nn3997), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3916), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_10|SUM_net ) );
      defparam ii3997.CONFIG_DATA = 16'h9A95;
      defparam ii3997.PLACE_LOCATION = "NONE";
      defparam ii3997.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3998 ( .DX(nn3998), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3917), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_11|SUM_net ) );
      defparam ii3998.CONFIG_DATA = 16'h9A95;
      defparam ii3998.PLACE_LOCATION = "NONE";
      defparam ii3998.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3999 ( .DX(nn3999), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3918), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_12|SUM_net ) );
      defparam ii3999.CONFIG_DATA = 16'h9A95;
      defparam ii3999.PLACE_LOCATION = "NONE";
      defparam ii3999.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4000 ( .DX(nn4000), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3919), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_13|SUM_net ) );
      defparam ii4000.CONFIG_DATA = 16'h9A95;
      defparam ii4000.PLACE_LOCATION = "NONE";
      defparam ii4000.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4001 ( .DX(nn4001), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn3920), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_14|SUM_net ) );
      defparam ii4001.CONFIG_DATA = 16'h9A95;
      defparam ii4001.PLACE_LOCATION = "NONE";
      defparam ii4001.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4002 ( .DX(nn4002), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(nn3868), .F2(dummy_488_), .F3(\coefcal1_divide_inst1_u116_XORCI_15|SUM_net ) );
      defparam ii4002.CONFIG_DATA = 16'h9A95;
      defparam ii4002.PLACE_LOCATION = "NONE";
      defparam ii4002.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4003 ( .DX(nn4003), .F0(dummy_abc_2674_), .F1(dummy_abc_2675_), .F2(dummy_abc_2676_), .F3(dummy_abc_2677_) );
      defparam ii4003.CONFIG_DATA = 16'hFFFF;
      defparam ii4003.PLACE_LOCATION = "NONE";
      defparam ii4003.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_39_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_507_ ), 
        .DX( {nn4003, nn4002, nn4001, nn4000, nn3999, nn3998, nn3997, nn3996, 
              nn3995, nn3994, nn3993, nn3992, nn3991, nn3990, nn3989, nn3988, 
              nn3987, nn3986} ), 
        .SUM( {\coefcal1_divide_inst1_u150_XORCI_17|SUM_net , dummy_508_, 
              dummy_509_, dummy_510_, dummy_511_, dummy_512_, dummy_513_, dummy_514_, 
              dummy_515_, dummy_516_, dummy_517_, dummy_518_, dummy_519_, dummy_520_, 
              dummy_521_, dummy_522_, dummy_523_, dummy_524_} )
      );
    CS_LUT4_PRIM ii4024 ( .DX(nn4024), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(dummy_507_), .F2(nn3984), .F3(dummy_abc_2678_) );
      defparam ii4024.CONFIG_DATA = 16'h5C5C;
      defparam ii4024.PLACE_LOCATION = "NONE";
      defparam ii4024.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4025 ( .DX(nn4025), .F0(rst), .F1(dummy_203_), .F2(nn3985), .F3(nn4024) );
      defparam ii4025.CONFIG_DATA = 16'hFFFB;
      defparam ii4025.PLACE_LOCATION = "NONE";
      defparam ii4025.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4026 ( .DX(nn4026), .F0(\cal1_u__reg[0]|Q_net ), .F1(nn4025), .F2(dummy_abc_2679_), .F3(dummy_abc_2680_) );
      defparam ii4026.CONFIG_DATA = 16'h6666;
      defparam ii4026.PLACE_LOCATION = "NONE";
      defparam ii4026.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4027 ( .DX(nn4027), .F0(rst), .F1(dummy_203_), .F2(nn3985), .F3(nn4024) );
      defparam ii4027.CONFIG_DATA = 16'hFFFB;
      defparam ii4027.PLACE_LOCATION = "NONE";
      defparam ii4027.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4028 ( .DX(nn4028), .F0(rst), .F1(\coefcal1_xDividend__reg[1]|Q_net ), .F2(\coefcal1_xDivisor__reg[0]|Q_net ), .F3(nn3984) );
      defparam ii4028.CONFIG_DATA = 16'h4055;
      defparam ii4028.PLACE_LOCATION = "NONE";
      defparam ii4028.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4029 ( .DX(nn4029), .F0(dummy_488_), .F1(dummy_203_), .F2(nn3984), .F3(nn4028) );
      defparam ii4029.CONFIG_DATA = 16'hC400;
      defparam ii4029.PLACE_LOCATION = "NONE";
      defparam ii4029.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4030 ( .DX(nn4030), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(dummy_469_), .F2(nn3984), .F3(dummy_abc_2681_) );
      defparam ii4030.CONFIG_DATA = 16'h5C5C;
      defparam ii4030.PLACE_LOCATION = "NONE";
      defparam ii4030.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4031 ( .DX(nn4031), .F0(rst), .F1(dummy_203_), .F2(nn3985), .F3(nn4030) );
      defparam ii4031.CONFIG_DATA = 16'h0004;
      defparam ii4031.PLACE_LOCATION = "NONE";
      defparam ii4031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4032 ( .DX(nn4032), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_450_), .F3(nn3984) );
      defparam ii4032.CONFIG_DATA = 16'h77F0;
      defparam ii4032.PLACE_LOCATION = "NONE";
      defparam ii4032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4033 ( .DX(nn4033), .F0(rst), .F1(dummy_203_), .F2(nn4032), .F3(dummy_abc_2682_) );
      defparam ii4033.CONFIG_DATA = 16'h0404;
      defparam ii4033.PLACE_LOCATION = "NONE";
      defparam ii4033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4034 ( .DX(nn4034), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(dummy_431_), .F2(nn3984), .F3(dummy_abc_2683_) );
      defparam ii4034.CONFIG_DATA = 16'h5C5C;
      defparam ii4034.PLACE_LOCATION = "NONE";
      defparam ii4034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4035 ( .DX(nn4035), .F0(rst), .F1(dummy_203_), .F2(nn3985), .F3(nn4034) );
      defparam ii4035.CONFIG_DATA = 16'h0004;
      defparam ii4035.PLACE_LOCATION = "NONE";
      defparam ii4035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4036 ( .DX(nn4036), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(dummy_412_), .F2(nn3984), .F3(dummy_abc_2684_) );
      defparam ii4036.CONFIG_DATA = 16'h5C5C;
      defparam ii4036.PLACE_LOCATION = "NONE";
      defparam ii4036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4037 ( .DX(nn4037), .F0(rst), .F1(dummy_203_), .F2(nn3985), .F3(nn4036) );
      defparam ii4037.CONFIG_DATA = 16'h0004;
      defparam ii4037.PLACE_LOCATION = "NONE";
      defparam ii4037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4038 ( .DX(nn4038), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_393_), .F3(nn3984) );
      defparam ii4038.CONFIG_DATA = 16'h880F;
      defparam ii4038.PLACE_LOCATION = "NONE";
      defparam ii4038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4039 ( .DX(nn4039), .F0(rst), .F1(dummy_203_), .F2(nn4038), .F3(dummy_abc_2685_) );
      defparam ii4039.CONFIG_DATA = 16'h4040;
      defparam ii4039.PLACE_LOCATION = "NONE";
      defparam ii4039.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4040 ( .DX(nn4040), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_374_), .F3(nn3984) );
      defparam ii4040.CONFIG_DATA = 16'h77F0;
      defparam ii4040.PLACE_LOCATION = "NONE";
      defparam ii4040.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4041 ( .DX(nn4041), .F0(rst), .F1(dummy_203_), .F2(nn4040), .F3(dummy_abc_2686_) );
      defparam ii4041.CONFIG_DATA = 16'h0404;
      defparam ii4041.PLACE_LOCATION = "NONE";
      defparam ii4041.PCK_LOCATION = "NONE";
    scaler_ipc_adder_8 carry_8 ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_dinxy_cen_cal1_u134_mac} ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_886_ ), 
        .DX( {nn4041, nn4039, nn4037, nn4035, nn4033, nn4031, nn4029, nn4027} ), 
        .SUM( {\coefcal1_u61_XORCI_7|SUM_net , \coefcal1_u61_XORCI_6|SUM_net , 
              \coefcal1_u61_XORCI_5|SUM_net , \coefcal1_u61_XORCI_4|SUM_net , 
              \coefcal1_u61_XORCI_3|SUM_net , \coefcal1_u61_XORCI_2|SUM_net , 
              \coefcal1_u61_XORCI_1|SUM_net , \coefcal1_u61_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4052 ( .DX(nn4052), .F0(\cal1_u__reg[1]|Q_net ), .F1(\coefcal1_u61_XORCI_1|SUM_net ), .F2(dummy_abc_2687_), .F3(dummy_abc_2688_) );
      defparam ii4052.CONFIG_DATA = 16'h6666;
      defparam ii4052.PLACE_LOCATION = "NONE";
      defparam ii4052.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4053 ( .DX(nn4053), .F0(\cal1_u__reg[2]|Q_net ), .F1(\coefcal1_u61_XORCI_2|SUM_net ), .F2(dummy_abc_2689_), .F3(dummy_abc_2690_) );
      defparam ii4053.CONFIG_DATA = 16'h6666;
      defparam ii4053.PLACE_LOCATION = "NONE";
      defparam ii4053.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4054 ( .DX(nn4054), .F0(\cal1_u__reg[3]|Q_net ), .F1(\coefcal1_u61_XORCI_3|SUM_net ), .F2(dummy_abc_2691_), .F3(dummy_abc_2692_) );
      defparam ii4054.CONFIG_DATA = 16'h6666;
      defparam ii4054.PLACE_LOCATION = "NONE";
      defparam ii4054.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4055 ( .DX(nn4055), .F0(\cal1_u__reg[4]|Q_net ), .F1(\coefcal1_u61_XORCI_4|SUM_net ), .F2(dummy_abc_2693_), .F3(dummy_abc_2694_) );
      defparam ii4055.CONFIG_DATA = 16'h6666;
      defparam ii4055.PLACE_LOCATION = "NONE";
      defparam ii4055.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4056 ( .DX(nn4056), .F0(\cal1_u__reg[5]|Q_net ), .F1(\coefcal1_u61_XORCI_5|SUM_net ), .F2(dummy_abc_2695_), .F3(dummy_abc_2696_) );
      defparam ii4056.CONFIG_DATA = 16'h6666;
      defparam ii4056.PLACE_LOCATION = "NONE";
      defparam ii4056.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4057 ( .DX(nn4057), .F0(\cal1_u__reg[6]|Q_net ), .F1(\coefcal1_u61_XORCI_6|SUM_net ), .F2(dummy_abc_2697_), .F3(dummy_abc_2698_) );
      defparam ii4057.CONFIG_DATA = 16'h6666;
      defparam ii4057.PLACE_LOCATION = "NONE";
      defparam ii4057.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4058 ( .DX(nn4058), .F0(\cal1_u__reg[7]|Q_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_abc_2699_), .F3(dummy_abc_2700_) );
      defparam ii4058.CONFIG_DATA = 16'h6666;
      defparam ii4058.PLACE_LOCATION = "NONE";
      defparam ii4058.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4059 ( .DX(nn4059), .F0(\cal1_u__reg[8]|Q_net ), .F1(dummy_abc_2701_), .F2(dummy_abc_2702_), .F3(dummy_abc_2703_) );
      defparam ii4059.CONFIG_DATA = 16'hAAAA;
      defparam ii4059.PLACE_LOCATION = "NONE";
      defparam ii4059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4060 ( .DX(nn4060), .F0(\cal1_u__reg[9]|Q_net ), .F1(dummy_abc_2704_), .F2(dummy_abc_2705_), .F3(dummy_abc_2706_) );
      defparam ii4060.CONFIG_DATA = 16'hAAAA;
      defparam ii4060.PLACE_LOCATION = "NONE";
      defparam ii4060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4061 ( .DX(nn4061), .F0(\cal1_u__reg[10]|Q_net ), .F1(dummy_abc_2707_), .F2(dummy_abc_2708_), .F3(dummy_abc_2709_) );
      defparam ii4061.CONFIG_DATA = 16'hAAAA;
      defparam ii4061.PLACE_LOCATION = "NONE";
      defparam ii4061.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4062 ( .DX(nn4062), .F0(\cal1_u__reg[11]|Q_net ), .F1(dummy_abc_2710_), .F2(dummy_abc_2711_), .F3(dummy_abc_2712_) );
      defparam ii4062.CONFIG_DATA = 16'hAAAA;
      defparam ii4062.PLACE_LOCATION = "NONE";
      defparam ii4062.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4063 ( .DX(nn4063), .F0(\cal1_u__reg[12]|Q_net ), .F1(dummy_abc_2713_), .F2(dummy_abc_2714_), .F3(dummy_abc_2715_) );
      defparam ii4063.CONFIG_DATA = 16'hAAAA;
      defparam ii4063.PLACE_LOCATION = "NONE";
      defparam ii4063.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4064 ( .DX(nn4064), .F0(\cal1_u__reg[13]|Q_net ), .F1(dummy_abc_2716_), .F2(dummy_abc_2717_), .F3(dummy_abc_2718_) );
      defparam ii4064.CONFIG_DATA = 16'hAAAA;
      defparam ii4064.PLACE_LOCATION = "NONE";
      defparam ii4064.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4065 ( .DX(nn4065), .F0(\cal1_u__reg[14]|Q_net ), .F1(dummy_abc_2719_), .F2(dummy_abc_2720_), .F3(dummy_abc_2721_) );
      defparam ii4065.CONFIG_DATA = 16'hAAAA;
      defparam ii4065.PLACE_LOCATION = "NONE";
      defparam ii4065.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4066 ( .DX(nn4066), .F0(\cal1_u__reg[15]|Q_net ), .F1(dummy_abc_2722_), .F2(dummy_abc_2723_), .F3(dummy_abc_2724_) );
      defparam ii4066.CONFIG_DATA = 16'hAAAA;
      defparam ii4066.PLACE_LOCATION = "NONE";
      defparam ii4066.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4067 ( .DX(nn4067), .F0(\cal1_u__reg[16]|Q_net ), .F1(dummy_abc_2725_), .F2(dummy_abc_2726_), .F3(dummy_abc_2727_) );
      defparam ii4067.CONFIG_DATA = 16'hAAAA;
      defparam ii4067.PLACE_LOCATION = "NONE";
      defparam ii4067.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17 ( 
        .CA( {\cal1_u__reg[16]|Q_net , \cal1_u__reg[15]|Q_net , 
              \cal1_u__reg[14]|Q_net , \cal1_u__reg[13]|Q_net , \cal1_u__reg[12]|Q_net , 
              \cal1_u__reg[11]|Q_net , \cal1_u__reg[10]|Q_net , \cal1_u__reg[9]|Q_net , 
              \cal1_u__reg[8]|Q_net , \cal1_u__reg[7]|Q_net , \cal1_u__reg[6]|Q_net , 
              \cal1_u__reg[5]|Q_net , \cal1_u__reg[4]|Q_net , \cal1_u__reg[3]|Q_net , 
              \cal1_u__reg[2]|Q_net , \cal1_u__reg[1]|Q_net , \cal1_u__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_138_ ), 
        .DX( {nn4067, nn4066, nn4065, nn4064, nn4063, nn4062, nn4061, nn4060, 
              nn4059, nn4058, nn4057, nn4056, nn4055, nn4054, nn4053, nn4052, 
              nn4026} ), 
        .SUM( {\cal1_u127_XORCI_16|SUM_net , \cal1_u127_XORCI_15|SUM_net , 
              \cal1_u127_XORCI_14|SUM_net , \cal1_u127_XORCI_13|SUM_net , \cal1_u127_XORCI_12|SUM_net , 
              \cal1_u127_XORCI_11|SUM_net , \cal1_u127_XORCI_10|SUM_net , \cal1_u127_XORCI_9|SUM_net , 
              \cal1_u127_XORCI_8|SUM_net , \cal1_u127_XORCI_7|SUM_net , \cal1_u127_XORCI_6|SUM_net , 
              \cal1_u127_XORCI_5|SUM_net , \cal1_u127_XORCI_4|SUM_net , \cal1_u127_XORCI_3|SUM_net , 
              \cal1_u127_XORCI_2|SUM_net , \cal1_u127_XORCI_1|SUM_net , \cal1_u127_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4087 ( .DX(nn4087), .F0(\cal1_u__reg[6]|Q_net ), .F1(\cal1_u__reg[7]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(\cal1_u127_XORCI_7|SUM_net ) );
      defparam ii4087.CONFIG_DATA = 16'hC639;
      defparam ii4087.PLACE_LOCATION = "NONE";
      defparam ii4087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4088 ( .DX(nn4088), .F0(\cal1_u__reg[6]|Q_net ), .F1(\cal1_u__reg[7]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(\cal1_u127_XORCI_7|SUM_net ) );
      defparam ii4088.CONFIG_DATA = 16'h08CE;
      defparam ii4088.PLACE_LOCATION = "NONE";
      defparam ii4088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4089 ( .DX(nn4089), .F0(\cal1_u__reg[8]|Q_net ), .F1(\cal1_u127_XORCI_8|SUM_net ), .F2(nn4087), .F3(nn4088) );
      defparam ii4089.CONFIG_DATA = 16'h6090;
      defparam ii4089.PLACE_LOCATION = "NONE";
      defparam ii4089.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4090 ( .DX(nn4090), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\cal1_u__reg[6]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(nn4089) );
      defparam ii4090.CONFIG_DATA = 16'h96AA;
      defparam ii4090.PLACE_LOCATION = "NONE";
      defparam ii4090.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4091 ( .DX(nn4091), .F0(dummy_35_), .F1(dummy_22_), .F2(nn4090), .F3(dummy_abc_2728_) );
      defparam ii4091.CONFIG_DATA = 16'h8080;
      defparam ii4091.PLACE_LOCATION = "NONE";
      defparam ii4091.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4092 ( .DX(nn4092), .F0(dummy_35_), .F1(dummy_22_), .F2(nn1312), .F3(dummy_abc_2729_) );
      defparam ii4092.CONFIG_DATA = 16'hF7F7;
      defparam ii4092.PLACE_LOCATION = "NONE";
      defparam ii4092.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4093 ( .DX(nn4093), .F0(dummy_52_), .F1(nn1329), .F2(nn4092), .F3(dummy_abc_2730_) );
      defparam ii4093.CONFIG_DATA = 16'hD0D0;
      defparam ii4093.PLACE_LOCATION = "NONE";
      defparam ii4093.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4094 ( .DX(nn4094), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\cal1_u__reg[6]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(nn4089) );
      defparam ii4094.CONFIG_DATA = 16'h96AA;
      defparam ii4094.PLACE_LOCATION = "NONE";
      defparam ii4094.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4095 ( .DX(nn4095), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(nn4089), .F2(dummy_abc_2731_), .F3(dummy_abc_2732_) );
      defparam ii4095.CONFIG_DATA = 16'h9999;
      defparam ii4095.PLACE_LOCATION = "NONE";
      defparam ii4095.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4096 ( .DX(nn4096), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(dummy_abc_2733_), .F2(dummy_abc_2734_), .F3(dummy_abc_2735_) );
      defparam ii4096.CONFIG_DATA = 16'hAAAA;
      defparam ii4096.PLACE_LOCATION = "NONE";
      defparam ii4096.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4097 ( .DX(nn4097), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(dummy_abc_2736_), .F2(dummy_abc_2737_), .F3(dummy_abc_2738_) );
      defparam ii4097.CONFIG_DATA = 16'hAAAA;
      defparam ii4097.PLACE_LOCATION = "NONE";
      defparam ii4097.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4098 ( .DX(nn4098), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(dummy_abc_2739_), .F2(dummy_abc_2740_), .F3(dummy_abc_2741_) );
      defparam ii4098.CONFIG_DATA = 16'hAAAA;
      defparam ii4098.PLACE_LOCATION = "NONE";
      defparam ii4098.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4099 ( .DX(nn4099), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(dummy_abc_2742_), .F2(dummy_abc_2743_), .F3(dummy_abc_2744_) );
      defparam ii4099.CONFIG_DATA = 16'hAAAA;
      defparam ii4099.PLACE_LOCATION = "NONE";
      defparam ii4099.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4100 ( .DX(nn4100), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(dummy_abc_2745_), .F2(dummy_abc_2746_), .F3(dummy_abc_2747_) );
      defparam ii4100.CONFIG_DATA = 16'hAAAA;
      defparam ii4100.PLACE_LOCATION = "NONE";
      defparam ii4100.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4101 ( .DX(nn4101), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(dummy_abc_2748_), .F2(dummy_abc_2749_), .F3(dummy_abc_2750_) );
      defparam ii4101.CONFIG_DATA = 16'hAAAA;
      defparam ii4101.PLACE_LOCATION = "NONE";
      defparam ii4101.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4102 ( .DX(nn4102), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(dummy_abc_2751_), .F2(dummy_abc_2752_), .F3(dummy_abc_2753_) );
      defparam ii4102.CONFIG_DATA = 16'hAAAA;
      defparam ii4102.PLACE_LOCATION = "NONE";
      defparam ii4102.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4103 ( .DX(nn4103), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(dummy_abc_2754_), .F2(dummy_abc_2755_), .F3(dummy_abc_2756_) );
      defparam ii4103.CONFIG_DATA = 16'hAAAA;
      defparam ii4103.PLACE_LOCATION = "NONE";
      defparam ii4103.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4104 ( .DX(nn4104), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(dummy_abc_2757_), .F2(dummy_abc_2758_), .F3(dummy_abc_2759_) );
      defparam ii4104.CONFIG_DATA = 16'hAAAA;
      defparam ii4104.PLACE_LOCATION = "NONE";
      defparam ii4104.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_1_ ( 
        .CA( {\cal1_ramRdAddr__reg[10]|Q_net , \cal1_ramRdAddr__reg[9]|Q_net , 
              \cal1_ramRdAddr__reg[8]|Q_net , \cal1_ramRdAddr__reg[7]|Q_net , 
              \cal1_ramRdAddr__reg[6]|Q_net , \cal1_ramRdAddr__reg[5]|Q_net , 
              \cal1_ramRdAddr__reg[4]|Q_net , \cal1_ramRdAddr__reg[3]|Q_net , 
              \cal1_ramRdAddr__reg[2]|Q_net , \cal1_ramRdAddr__reg[1]|Q_net , 
              \cal1_ramRdAddr__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_13_ ), 
        .DX( {nn4104, nn4103, nn4102, nn4101, nn4100, nn4099, nn4098, nn4097, 
              nn4096, nn4095, nn4094} ), 
        .SUM( {\cal1_u130_XORCI_10|SUM_net , \cal1_u130_XORCI_9|SUM_net , 
              \cal1_u130_XORCI_8|SUM_net , \cal1_u130_XORCI_7|SUM_net , \cal1_u130_XORCI_6|SUM_net , 
              \cal1_u130_XORCI_5|SUM_net , \cal1_u130_XORCI_4|SUM_net , \cal1_u130_XORCI_3|SUM_net , 
              \cal1_u130_XORCI_2|SUM_net , \cal1_u130_XORCI_1|SUM_net , \cal1_u130_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4118 ( .DX(nn4118), .F0(\cal1_u130_XORCI_10|SUM_net ), .F1(nn1329), .F2(dummy_abc_2760_), .F3(dummy_abc_2761_) );
      defparam ii4118.CONFIG_DATA = 16'h2222;
      defparam ii4118.PLACE_LOCATION = "NONE";
      defparam ii4118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4119 ( .DX(nn4119), .F0(\cal1_u130_XORCI_1|SUM_net ), .F1(nn1329), .F2(dummy_abc_2762_), .F3(dummy_abc_2763_) );
      defparam ii4119.CONFIG_DATA = 16'h2222;
      defparam ii4119.PLACE_LOCATION = "NONE";
      defparam ii4119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4120 ( .DX(nn4120), .F0(\cal1_u130_XORCI_2|SUM_net ), .F1(nn1329), .F2(dummy_abc_2764_), .F3(dummy_abc_2765_) );
      defparam ii4120.CONFIG_DATA = 16'h2222;
      defparam ii4120.PLACE_LOCATION = "NONE";
      defparam ii4120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4121 ( .DX(nn4121), .F0(\cal1_u130_XORCI_3|SUM_net ), .F1(nn1329), .F2(dummy_abc_2766_), .F3(dummy_abc_2767_) );
      defparam ii4121.CONFIG_DATA = 16'h2222;
      defparam ii4121.PLACE_LOCATION = "NONE";
      defparam ii4121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4122 ( .DX(nn4122), .F0(\cal1_u130_XORCI_4|SUM_net ), .F1(nn1329), .F2(dummy_abc_2768_), .F3(dummy_abc_2769_) );
      defparam ii4122.CONFIG_DATA = 16'h2222;
      defparam ii4122.PLACE_LOCATION = "NONE";
      defparam ii4122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4123 ( .DX(nn4123), .F0(\cal1_u130_XORCI_5|SUM_net ), .F1(nn1329), .F2(dummy_abc_2770_), .F3(dummy_abc_2771_) );
      defparam ii4123.CONFIG_DATA = 16'h2222;
      defparam ii4123.PLACE_LOCATION = "NONE";
      defparam ii4123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4124 ( .DX(nn4124), .F0(\cal1_u130_XORCI_6|SUM_net ), .F1(nn1329), .F2(dummy_abc_2772_), .F3(dummy_abc_2773_) );
      defparam ii4124.CONFIG_DATA = 16'h2222;
      defparam ii4124.PLACE_LOCATION = "NONE";
      defparam ii4124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4125 ( .DX(nn4125), .F0(\cal1_u130_XORCI_7|SUM_net ), .F1(nn1329), .F2(dummy_abc_2774_), .F3(dummy_abc_2775_) );
      defparam ii4125.CONFIG_DATA = 16'h2222;
      defparam ii4125.PLACE_LOCATION = "NONE";
      defparam ii4125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4126 ( .DX(nn4126), .F0(\cal1_u130_XORCI_8|SUM_net ), .F1(nn1329), .F2(dummy_abc_2776_), .F3(dummy_abc_2777_) );
      defparam ii4126.CONFIG_DATA = 16'h2222;
      defparam ii4126.PLACE_LOCATION = "NONE";
      defparam ii4126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4127 ( .DX(nn4127), .F0(\cal1_u130_XORCI_9|SUM_net ), .F1(nn1329), .F2(dummy_abc_2778_), .F3(dummy_abc_2779_) );
      defparam ii4127.CONFIG_DATA = 16'h2222;
      defparam ii4127.PLACE_LOCATION = "NONE";
      defparam ii4127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4128 ( .DX(nn4128), .F0(\cal1_u__reg[0]|Q_net ), .F1(nn4025), .F2(dummy_abc_2780_), .F3(dummy_abc_2781_) );
      defparam ii4128.CONFIG_DATA = 16'h6666;
      defparam ii4128.PLACE_LOCATION = "NONE";
      defparam ii4128.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4129 ( .DX(nn4129), .F0(nn4128), .F1(nn1329), .F2(dummy_abc_2782_), .F3(dummy_abc_2783_) );
      defparam ii4129.CONFIG_DATA = 16'h2222;
      defparam ii4129.PLACE_LOCATION = "NONE";
      defparam ii4129.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4130 ( .DX(nn4130), .F0(\cal1_u127_XORCI_10|SUM_net ), .F1(nn1329), .F2(dummy_abc_2784_), .F3(dummy_abc_2785_) );
      defparam ii4130.CONFIG_DATA = 16'h2222;
      defparam ii4130.PLACE_LOCATION = "NONE";
      defparam ii4130.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4131 ( .DX(nn4131), .F0(\cal1_u127_XORCI_11|SUM_net ), .F1(nn1329), .F2(dummy_abc_2786_), .F3(dummy_abc_2787_) );
      defparam ii4131.CONFIG_DATA = 16'h2222;
      defparam ii4131.PLACE_LOCATION = "NONE";
      defparam ii4131.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4132 ( .DX(nn4132), .F0(\cal1_u127_XORCI_12|SUM_net ), .F1(nn1329), .F2(dummy_abc_2788_), .F3(dummy_abc_2789_) );
      defparam ii4132.CONFIG_DATA = 16'h2222;
      defparam ii4132.PLACE_LOCATION = "NONE";
      defparam ii4132.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4133 ( .DX(nn4133), .F0(\cal1_u127_XORCI_13|SUM_net ), .F1(nn1329), .F2(dummy_abc_2790_), .F3(dummy_abc_2791_) );
      defparam ii4133.CONFIG_DATA = 16'h2222;
      defparam ii4133.PLACE_LOCATION = "NONE";
      defparam ii4133.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4134 ( .DX(nn4134), .F0(\cal1_u127_XORCI_14|SUM_net ), .F1(nn1329), .F2(dummy_abc_2792_), .F3(dummy_abc_2793_) );
      defparam ii4134.CONFIG_DATA = 16'h2222;
      defparam ii4134.PLACE_LOCATION = "NONE";
      defparam ii4134.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4135 ( .DX(nn4135), .F0(\cal1_u127_XORCI_15|SUM_net ), .F1(nn1329), .F2(dummy_abc_2794_), .F3(dummy_abc_2795_) );
      defparam ii4135.CONFIG_DATA = 16'h2222;
      defparam ii4135.PLACE_LOCATION = "NONE";
      defparam ii4135.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4136 ( .DX(nn4136), .F0(\cal1_u127_XORCI_16|SUM_net ), .F1(nn1329), .F2(dummy_abc_2796_), .F3(dummy_abc_2797_) );
      defparam ii4136.CONFIG_DATA = 16'h2222;
      defparam ii4136.PLACE_LOCATION = "NONE";
      defparam ii4136.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4137 ( .DX(nn4137), .F0(\cal1_u127_XORCI_1|SUM_net ), .F1(nn1329), .F2(dummy_abc_2798_), .F3(dummy_abc_2799_) );
      defparam ii4137.CONFIG_DATA = 16'h2222;
      defparam ii4137.PLACE_LOCATION = "NONE";
      defparam ii4137.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4138 ( .DX(nn4138), .F0(\cal1_u127_XORCI_2|SUM_net ), .F1(nn1329), .F2(dummy_abc_2800_), .F3(dummy_abc_2801_) );
      defparam ii4138.CONFIG_DATA = 16'h2222;
      defparam ii4138.PLACE_LOCATION = "NONE";
      defparam ii4138.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4139 ( .DX(nn4139), .F0(\cal1_u127_XORCI_3|SUM_net ), .F1(nn1329), .F2(dummy_abc_2802_), .F3(dummy_abc_2803_) );
      defparam ii4139.CONFIG_DATA = 16'h2222;
      defparam ii4139.PLACE_LOCATION = "NONE";
      defparam ii4139.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4140 ( .DX(nn4140), .F0(\cal1_u127_XORCI_4|SUM_net ), .F1(nn1329), .F2(dummy_abc_2804_), .F3(dummy_abc_2805_) );
      defparam ii4140.CONFIG_DATA = 16'h2222;
      defparam ii4140.PLACE_LOCATION = "NONE";
      defparam ii4140.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4141 ( .DX(nn4141), .F0(\cal1_u127_XORCI_5|SUM_net ), .F1(nn1329), .F2(dummy_abc_2806_), .F3(dummy_abc_2807_) );
      defparam ii4141.CONFIG_DATA = 16'h2222;
      defparam ii4141.PLACE_LOCATION = "NONE";
      defparam ii4141.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4142 ( .DX(nn4142), .F0(\cal1_u127_XORCI_6|SUM_net ), .F1(nn1329), .F2(dummy_abc_2808_), .F3(dummy_abc_2809_) );
      defparam ii4142.CONFIG_DATA = 16'h2222;
      defparam ii4142.PLACE_LOCATION = "NONE";
      defparam ii4142.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4143 ( .DX(nn4143), .F0(\cal1_u127_XORCI_7|SUM_net ), .F1(nn1329), .F2(dummy_abc_2810_), .F3(dummy_abc_2811_) );
      defparam ii4143.CONFIG_DATA = 16'h2222;
      defparam ii4143.PLACE_LOCATION = "NONE";
      defparam ii4143.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4144 ( .DX(nn4144), .F0(\cal1_u127_XORCI_8|SUM_net ), .F1(nn1329), .F2(dummy_abc_2812_), .F3(dummy_abc_2813_) );
      defparam ii4144.CONFIG_DATA = 16'h2222;
      defparam ii4144.PLACE_LOCATION = "NONE";
      defparam ii4144.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4145 ( .DX(nn4145), .F0(\cal1_u127_XORCI_9|SUM_net ), .F1(nn1329), .F2(dummy_abc_2814_), .F3(dummy_abc_2815_) );
      defparam ii4145.CONFIG_DATA = 16'h2222;
      defparam ii4145.PLACE_LOCATION = "NONE";
      defparam ii4145.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4146 ( .DX(nn4146), .F0(rst), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_526_), .F3(nn2644) );
      defparam ii4146.CONFIG_DATA = 16'h3363;
      defparam ii4146.PLACE_LOCATION = "NONE";
      defparam ii4146.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4147 ( .DX(nn4147), .F0(dummy_35_), .F1(nn4146), .F2(dummy_abc_2816_), .F3(dummy_abc_2817_) );
      defparam ii4147.CONFIG_DATA = 16'h8888;
      defparam ii4147.PLACE_LOCATION = "NONE";
      defparam ii4147.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4148 ( .DX(nn4148), .F0(dummy_35_), .F1(\cal1_u128_XORCI_10|SUM_net ), .F2(dummy_abc_2818_), .F3(dummy_abc_2819_) );
      defparam ii4148.CONFIG_DATA = 16'h8888;
      defparam ii4148.PLACE_LOCATION = "NONE";
      defparam ii4148.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4149 ( .DX(nn4149), .F0(dummy_35_), .F1(\cal1_u128_XORCI_11|SUM_net ), .F2(dummy_abc_2820_), .F3(dummy_abc_2821_) );
      defparam ii4149.CONFIG_DATA = 16'h8888;
      defparam ii4149.PLACE_LOCATION = "NONE";
      defparam ii4149.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4150 ( .DX(nn4150), .F0(dummy_35_), .F1(\cal1_u128_XORCI_12|SUM_net ), .F2(dummy_abc_2822_), .F3(dummy_abc_2823_) );
      defparam ii4150.CONFIG_DATA = 16'h8888;
      defparam ii4150.PLACE_LOCATION = "NONE";
      defparam ii4150.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4151 ( .DX(nn4151), .F0(dummy_35_), .F1(\cal1_u128_XORCI_13|SUM_net ), .F2(dummy_abc_2824_), .F3(dummy_abc_2825_) );
      defparam ii4151.CONFIG_DATA = 16'h8888;
      defparam ii4151.PLACE_LOCATION = "NONE";
      defparam ii4151.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4152 ( .DX(nn4152), .F0(dummy_35_), .F1(\cal1_u128_XORCI_14|SUM_net ), .F2(dummy_abc_2826_), .F3(dummy_abc_2827_) );
      defparam ii4152.CONFIG_DATA = 16'h8888;
      defparam ii4152.PLACE_LOCATION = "NONE";
      defparam ii4152.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4153 ( .DX(nn4153), .F0(dummy_35_), .F1(\cal1_u128_XORCI_15|SUM_net ), .F2(dummy_abc_2828_), .F3(dummy_abc_2829_) );
      defparam ii4153.CONFIG_DATA = 16'h8888;
      defparam ii4153.PLACE_LOCATION = "NONE";
      defparam ii4153.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4154 ( .DX(nn4154), .F0(dummy_35_), .F1(\cal1_u128_XORCI_16|SUM_net ), .F2(dummy_abc_2830_), .F3(dummy_abc_2831_) );
      defparam ii4154.CONFIG_DATA = 16'h8888;
      defparam ii4154.PLACE_LOCATION = "NONE";
      defparam ii4154.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4155 ( .DX(nn4155), .F0(dummy_35_), .F1(\cal1_u128_XORCI_1|SUM_net ), .F2(dummy_abc_2832_), .F3(dummy_abc_2833_) );
      defparam ii4155.CONFIG_DATA = 16'h8888;
      defparam ii4155.PLACE_LOCATION = "NONE";
      defparam ii4155.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4156 ( .DX(nn4156), .F0(dummy_35_), .F1(\cal1_u128_XORCI_2|SUM_net ), .F2(dummy_abc_2834_), .F3(dummy_abc_2835_) );
      defparam ii4156.CONFIG_DATA = 16'h8888;
      defparam ii4156.PLACE_LOCATION = "NONE";
      defparam ii4156.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4157 ( .DX(nn4157), .F0(dummy_35_), .F1(\cal1_u128_XORCI_3|SUM_net ), .F2(dummy_abc_2836_), .F3(dummy_abc_2837_) );
      defparam ii4157.CONFIG_DATA = 16'h8888;
      defparam ii4157.PLACE_LOCATION = "NONE";
      defparam ii4157.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4158 ( .DX(nn4158), .F0(dummy_35_), .F1(\cal1_u128_XORCI_4|SUM_net ), .F2(dummy_abc_2838_), .F3(dummy_abc_2839_) );
      defparam ii4158.CONFIG_DATA = 16'h8888;
      defparam ii4158.PLACE_LOCATION = "NONE";
      defparam ii4158.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4159 ( .DX(nn4159), .F0(dummy_35_), .F1(\cal1_u128_XORCI_5|SUM_net ), .F2(dummy_abc_2840_), .F3(dummy_abc_2841_) );
      defparam ii4159.CONFIG_DATA = 16'h8888;
      defparam ii4159.PLACE_LOCATION = "NONE";
      defparam ii4159.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4160 ( .DX(nn4160), .F0(dummy_35_), .F1(\cal1_u128_XORCI_6|SUM_net ), .F2(dummy_abc_2842_), .F3(dummy_abc_2843_) );
      defparam ii4160.CONFIG_DATA = 16'h8888;
      defparam ii4160.PLACE_LOCATION = "NONE";
      defparam ii4160.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4161 ( .DX(nn4161), .F0(dummy_35_), .F1(\cal1_u128_XORCI_7|SUM_net ), .F2(dummy_abc_2844_), .F3(dummy_abc_2845_) );
      defparam ii4161.CONFIG_DATA = 16'h8888;
      defparam ii4161.PLACE_LOCATION = "NONE";
      defparam ii4161.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4162 ( .DX(nn4162), .F0(dummy_35_), .F1(\cal1_u128_XORCI_8|SUM_net ), .F2(dummy_abc_2846_), .F3(dummy_abc_2847_) );
      defparam ii4162.CONFIG_DATA = 16'h8888;
      defparam ii4162.PLACE_LOCATION = "NONE";
      defparam ii4162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4163 ( .DX(nn4163), .F0(dummy_35_), .F1(\cal1_u128_XORCI_9|SUM_net ), .F2(dummy_abc_2848_), .F3(dummy_abc_2849_) );
      defparam ii4163.CONFIG_DATA = 16'h8888;
      defparam ii4163.PLACE_LOCATION = "NONE";
      defparam ii4163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4164 ( .DX(nn4164), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(nn1329), .F2(dummy_abc_2850_), .F3(dummy_abc_2851_) );
      defparam ii4164.CONFIG_DATA = 16'h1111;
      defparam ii4164.PLACE_LOCATION = "NONE";
      defparam ii4164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4165 ( .DX(nn4165), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_2852_), .F2(dummy_abc_2853_), .F3(dummy_abc_2854_) );
      defparam ii4165.CONFIG_DATA = 16'h5555;
      defparam ii4165.PLACE_LOCATION = "NONE";
      defparam ii4165.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4166 ( .DX(nn4166), .F0(\cal1_xAddress__reg[1]|Q_net ), .F1(dummy_abc_2855_), .F2(dummy_abc_2856_), .F3(dummy_abc_2857_) );
      defparam ii4166.CONFIG_DATA = 16'hAAAA;
      defparam ii4166.PLACE_LOCATION = "NONE";
      defparam ii4166.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4167 ( .DX(nn4167), .F0(\cal1_xAddress__reg[2]|Q_net ), .F1(dummy_abc_2858_), .F2(dummy_abc_2859_), .F3(dummy_abc_2860_) );
      defparam ii4167.CONFIG_DATA = 16'hAAAA;
      defparam ii4167.PLACE_LOCATION = "NONE";
      defparam ii4167.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4168 ( .DX(nn4168), .F0(\cal1_xAddress__reg[3]|Q_net ), .F1(dummy_abc_2861_), .F2(dummy_abc_2862_), .F3(dummy_abc_2863_) );
      defparam ii4168.CONFIG_DATA = 16'hAAAA;
      defparam ii4168.PLACE_LOCATION = "NONE";
      defparam ii4168.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4169 ( .DX(nn4169), .F0(\cal1_xAddress__reg[4]|Q_net ), .F1(dummy_abc_2864_), .F2(dummy_abc_2865_), .F3(dummy_abc_2866_) );
      defparam ii4169.CONFIG_DATA = 16'hAAAA;
      defparam ii4169.PLACE_LOCATION = "NONE";
      defparam ii4169.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4170 ( .DX(nn4170), .F0(\cal1_xAddress__reg[5]|Q_net ), .F1(dummy_abc_2867_), .F2(dummy_abc_2868_), .F3(dummy_abc_2869_) );
      defparam ii4170.CONFIG_DATA = 16'hAAAA;
      defparam ii4170.PLACE_LOCATION = "NONE";
      defparam ii4170.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4171 ( .DX(nn4171), .F0(\cal1_xAddress__reg[6]|Q_net ), .F1(dummy_abc_2870_), .F2(dummy_abc_2871_), .F3(dummy_abc_2872_) );
      defparam ii4171.CONFIG_DATA = 16'hAAAA;
      defparam ii4171.PLACE_LOCATION = "NONE";
      defparam ii4171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4172 ( .DX(nn4172), .F0(\cal1_xAddress__reg[7]|Q_net ), .F1(dummy_abc_2873_), .F2(dummy_abc_2874_), .F3(dummy_abc_2875_) );
      defparam ii4172.CONFIG_DATA = 16'hAAAA;
      defparam ii4172.PLACE_LOCATION = "NONE";
      defparam ii4172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4173 ( .DX(nn4173), .F0(\cal1_xAddress__reg[8]|Q_net ), .F1(dummy_abc_2876_), .F2(dummy_abc_2877_), .F3(dummy_abc_2878_) );
      defparam ii4173.CONFIG_DATA = 16'hAAAA;
      defparam ii4173.PLACE_LOCATION = "NONE";
      defparam ii4173.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4174 ( .DX(nn4174), .F0(\cal1_xAddress__reg[9]|Q_net ), .F1(dummy_abc_2879_), .F2(dummy_abc_2880_), .F3(dummy_abc_2881_) );
      defparam ii4174.CONFIG_DATA = 16'hAAAA;
      defparam ii4174.PLACE_LOCATION = "NONE";
      defparam ii4174.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4175 ( .DX(nn4175), .F0(\cal1_xAddress__reg[10]|Q_net ), .F1(dummy_abc_2882_), .F2(dummy_abc_2883_), .F3(dummy_abc_2884_) );
      defparam ii4175.CONFIG_DATA = 16'hAAAA;
      defparam ii4175.PLACE_LOCATION = "NONE";
      defparam ii4175.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_2_ ( 
        .CA( {\cal1_xAddress__reg[10]|Q_net , \cal1_xAddress__reg[9]|Q_net , 
              \cal1_xAddress__reg[8]|Q_net , \cal1_xAddress__reg[7]|Q_net , 
              \cal1_xAddress__reg[6]|Q_net , \cal1_xAddress__reg[5]|Q_net , 
              \cal1_xAddress__reg[4]|Q_net , \cal1_xAddress__reg[3]|Q_net , 
              \cal1_xAddress__reg[2]|Q_net , \cal1_xAddress__reg[1]|Q_net , 
              \cal1_xAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_14_ ), 
        .DX( {nn4175, nn4174, nn4173, nn4172, nn4171, nn4170, nn4169, nn4168, 
              nn4167, nn4166, nn4165} ), 
        .SUM( {\cal1_u131_XORCI_10|SUM_net , \cal1_u131_XORCI_9|SUM_net , 
              \cal1_u131_XORCI_8|SUM_net , \cal1_u131_XORCI_7|SUM_net , \cal1_u131_XORCI_6|SUM_net , 
              \cal1_u131_XORCI_5|SUM_net , \cal1_u131_XORCI_4|SUM_net , \cal1_u131_XORCI_3|SUM_net , 
              \cal1_u131_XORCI_2|SUM_net , \cal1_u131_XORCI_1|SUM_net , \cal1_u131_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4189 ( .DX(nn4189), .F0(\cal1_u131_XORCI_10|SUM_net ), .F1(nn1329), .F2(dummy_abc_2885_), .F3(dummy_abc_2886_) );
      defparam ii4189.CONFIG_DATA = 16'h2222;
      defparam ii4189.PLACE_LOCATION = "NONE";
      defparam ii4189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4190 ( .DX(nn4190), .F0(\cal1_u131_XORCI_1|SUM_net ), .F1(nn1329), .F2(dummy_abc_2887_), .F3(dummy_abc_2888_) );
      defparam ii4190.CONFIG_DATA = 16'h2222;
      defparam ii4190.PLACE_LOCATION = "NONE";
      defparam ii4190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4191 ( .DX(nn4191), .F0(\cal1_u131_XORCI_2|SUM_net ), .F1(nn1329), .F2(dummy_abc_2889_), .F3(dummy_abc_2890_) );
      defparam ii4191.CONFIG_DATA = 16'h2222;
      defparam ii4191.PLACE_LOCATION = "NONE";
      defparam ii4191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4192 ( .DX(nn4192), .F0(\cal1_u131_XORCI_3|SUM_net ), .F1(nn1329), .F2(dummy_abc_2891_), .F3(dummy_abc_2892_) );
      defparam ii4192.CONFIG_DATA = 16'h2222;
      defparam ii4192.PLACE_LOCATION = "NONE";
      defparam ii4192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4193 ( .DX(nn4193), .F0(\cal1_u131_XORCI_4|SUM_net ), .F1(nn1329), .F2(dummy_abc_2893_), .F3(dummy_abc_2894_) );
      defparam ii4193.CONFIG_DATA = 16'h2222;
      defparam ii4193.PLACE_LOCATION = "NONE";
      defparam ii4193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4194 ( .DX(nn4194), .F0(\cal1_u131_XORCI_5|SUM_net ), .F1(nn1329), .F2(dummy_abc_2895_), .F3(dummy_abc_2896_) );
      defparam ii4194.CONFIG_DATA = 16'h2222;
      defparam ii4194.PLACE_LOCATION = "NONE";
      defparam ii4194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4195 ( .DX(nn4195), .F0(\cal1_u131_XORCI_6|SUM_net ), .F1(nn1329), .F2(dummy_abc_2897_), .F3(dummy_abc_2898_) );
      defparam ii4195.CONFIG_DATA = 16'h2222;
      defparam ii4195.PLACE_LOCATION = "NONE";
      defparam ii4195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4196 ( .DX(nn4196), .F0(\cal1_u131_XORCI_7|SUM_net ), .F1(nn1329), .F2(dummy_abc_2899_), .F3(dummy_abc_2900_) );
      defparam ii4196.CONFIG_DATA = 16'h2222;
      defparam ii4196.PLACE_LOCATION = "NONE";
      defparam ii4196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4197 ( .DX(nn4197), .F0(\cal1_u131_XORCI_8|SUM_net ), .F1(nn1329), .F2(dummy_abc_2901_), .F3(dummy_abc_2902_) );
      defparam ii4197.CONFIG_DATA = 16'h2222;
      defparam ii4197.PLACE_LOCATION = "NONE";
      defparam ii4197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4198 ( .DX(nn4198), .F0(\cal1_u131_XORCI_9|SUM_net ), .F1(nn1329), .F2(dummy_abc_2903_), .F3(dummy_abc_2904_) );
      defparam ii4198.CONFIG_DATA = 16'h2222;
      defparam ii4198.PLACE_LOCATION = "NONE";
      defparam ii4198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4199 ( .DX(nn4199), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(dummy_35_), .F2(dummy_abc_2905_), .F3(dummy_abc_2906_) );
      defparam ii4199.CONFIG_DATA = 16'h7777;
      defparam ii4199.PLACE_LOCATION = "NONE";
      defparam ii4199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4200 ( .DX(nn4200), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_2907_), .F2(dummy_abc_2908_), .F3(dummy_abc_2909_) );
      defparam ii4200.CONFIG_DATA = 16'h5555;
      defparam ii4200.PLACE_LOCATION = "NONE";
      defparam ii4200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4201 ( .DX(nn4201), .F0(\cal1_yAddress__reg[1]|Q_net ), .F1(dummy_abc_2910_), .F2(dummy_abc_2911_), .F3(dummy_abc_2912_) );
      defparam ii4201.CONFIG_DATA = 16'hAAAA;
      defparam ii4201.PLACE_LOCATION = "NONE";
      defparam ii4201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4202 ( .DX(nn4202), .F0(\cal1_yAddress__reg[2]|Q_net ), .F1(dummy_abc_2913_), .F2(dummy_abc_2914_), .F3(dummy_abc_2915_) );
      defparam ii4202.CONFIG_DATA = 16'hAAAA;
      defparam ii4202.PLACE_LOCATION = "NONE";
      defparam ii4202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4203 ( .DX(nn4203), .F0(\cal1_yAddress__reg[3]|Q_net ), .F1(dummy_abc_2916_), .F2(dummy_abc_2917_), .F3(dummy_abc_2918_) );
      defparam ii4203.CONFIG_DATA = 16'hAAAA;
      defparam ii4203.PLACE_LOCATION = "NONE";
      defparam ii4203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4204 ( .DX(nn4204), .F0(\cal1_yAddress__reg[4]|Q_net ), .F1(dummy_abc_2919_), .F2(dummy_abc_2920_), .F3(dummy_abc_2921_) );
      defparam ii4204.CONFIG_DATA = 16'hAAAA;
      defparam ii4204.PLACE_LOCATION = "NONE";
      defparam ii4204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4205 ( .DX(nn4205), .F0(\cal1_yAddress__reg[5]|Q_net ), .F1(dummy_abc_2922_), .F2(dummy_abc_2923_), .F3(dummy_abc_2924_) );
      defparam ii4205.CONFIG_DATA = 16'hAAAA;
      defparam ii4205.PLACE_LOCATION = "NONE";
      defparam ii4205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4206 ( .DX(nn4206), .F0(\cal1_yAddress__reg[6]|Q_net ), .F1(dummy_abc_2925_), .F2(dummy_abc_2926_), .F3(dummy_abc_2927_) );
      defparam ii4206.CONFIG_DATA = 16'hAAAA;
      defparam ii4206.PLACE_LOCATION = "NONE";
      defparam ii4206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4207 ( .DX(nn4207), .F0(\cal1_yAddress__reg[7]|Q_net ), .F1(dummy_abc_2928_), .F2(dummy_abc_2929_), .F3(dummy_abc_2930_) );
      defparam ii4207.CONFIG_DATA = 16'hAAAA;
      defparam ii4207.PLACE_LOCATION = "NONE";
      defparam ii4207.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4208 ( .DX(nn4208), .F0(\cal1_yAddress__reg[8]|Q_net ), .F1(dummy_abc_2931_), .F2(dummy_abc_2932_), .F3(dummy_abc_2933_) );
      defparam ii4208.CONFIG_DATA = 16'hAAAA;
      defparam ii4208.PLACE_LOCATION = "NONE";
      defparam ii4208.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4209 ( .DX(nn4209), .F0(\cal1_yAddress__reg[9]|Q_net ), .F1(dummy_abc_2934_), .F2(dummy_abc_2935_), .F3(dummy_abc_2936_) );
      defparam ii4209.CONFIG_DATA = 16'hAAAA;
      defparam ii4209.PLACE_LOCATION = "NONE";
      defparam ii4209.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4210 ( .DX(nn4210), .F0(\cal1_yAddress__reg[10]|Q_net ), .F1(dummy_abc_2937_), .F2(dummy_abc_2938_), .F3(dummy_abc_2939_) );
      defparam ii4210.CONFIG_DATA = 16'hAAAA;
      defparam ii4210.PLACE_LOCATION = "NONE";
      defparam ii4210.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_3_ ( 
        .CA( {\cal1_yAddress__reg[10]|Q_net , \cal1_yAddress__reg[9]|Q_net , 
              \cal1_yAddress__reg[8]|Q_net , \cal1_yAddress__reg[7]|Q_net , 
              \cal1_yAddress__reg[6]|Q_net , \cal1_yAddress__reg[5]|Q_net , 
              \cal1_yAddress__reg[4]|Q_net , \cal1_yAddress__reg[3]|Q_net , 
              \cal1_yAddress__reg[2]|Q_net , \cal1_yAddress__reg[1]|Q_net , 
              \cal1_yAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_15_ ), 
        .DX( {nn4210, nn4209, nn4208, nn4207, nn4206, nn4205, nn4204, nn4203, 
              nn4202, nn4201, nn4200} ), 
        .SUM( {\cal1_u132_XORCI_10|SUM_net , \cal1_u132_XORCI_9|SUM_net , 
              \cal1_u132_XORCI_8|SUM_net , \cal1_u132_XORCI_7|SUM_net , \cal1_u132_XORCI_6|SUM_net , 
              \cal1_u132_XORCI_5|SUM_net , \cal1_u132_XORCI_4|SUM_net , \cal1_u132_XORCI_3|SUM_net , 
              \cal1_u132_XORCI_2|SUM_net , \cal1_u132_XORCI_1|SUM_net , \cal1_u132_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4224 ( .DX(nn4224), .F0(dummy_35_), .F1(\cal1_u132_XORCI_10|SUM_net ), .F2(dummy_abc_2940_), .F3(dummy_abc_2941_) );
      defparam ii4224.CONFIG_DATA = 16'h8888;
      defparam ii4224.PLACE_LOCATION = "NONE";
      defparam ii4224.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4225 ( .DX(nn4225), .F0(dummy_35_), .F1(\cal1_u132_XORCI_1|SUM_net ), .F2(dummy_abc_2942_), .F3(dummy_abc_2943_) );
      defparam ii4225.CONFIG_DATA = 16'h8888;
      defparam ii4225.PLACE_LOCATION = "NONE";
      defparam ii4225.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4226 ( .DX(nn4226), .F0(dummy_35_), .F1(\cal1_u132_XORCI_2|SUM_net ), .F2(dummy_abc_2944_), .F3(dummy_abc_2945_) );
      defparam ii4226.CONFIG_DATA = 16'h8888;
      defparam ii4226.PLACE_LOCATION = "NONE";
      defparam ii4226.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4227 ( .DX(nn4227), .F0(dummy_35_), .F1(\cal1_u132_XORCI_3|SUM_net ), .F2(dummy_abc_2946_), .F3(dummy_abc_2947_) );
      defparam ii4227.CONFIG_DATA = 16'h8888;
      defparam ii4227.PLACE_LOCATION = "NONE";
      defparam ii4227.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4228 ( .DX(nn4228), .F0(dummy_35_), .F1(\cal1_u132_XORCI_4|SUM_net ), .F2(dummy_abc_2948_), .F3(dummy_abc_2949_) );
      defparam ii4228.CONFIG_DATA = 16'h8888;
      defparam ii4228.PLACE_LOCATION = "NONE";
      defparam ii4228.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4229 ( .DX(nn4229), .F0(dummy_35_), .F1(\cal1_u132_XORCI_5|SUM_net ), .F2(dummy_abc_2950_), .F3(dummy_abc_2951_) );
      defparam ii4229.CONFIG_DATA = 16'h8888;
      defparam ii4229.PLACE_LOCATION = "NONE";
      defparam ii4229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4230 ( .DX(nn4230), .F0(dummy_35_), .F1(\cal1_u132_XORCI_6|SUM_net ), .F2(dummy_abc_2952_), .F3(dummy_abc_2953_) );
      defparam ii4230.CONFIG_DATA = 16'h8888;
      defparam ii4230.PLACE_LOCATION = "NONE";
      defparam ii4230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4231 ( .DX(nn4231), .F0(dummy_35_), .F1(\cal1_u132_XORCI_7|SUM_net ), .F2(dummy_abc_2954_), .F3(dummy_abc_2955_) );
      defparam ii4231.CONFIG_DATA = 16'h8888;
      defparam ii4231.PLACE_LOCATION = "NONE";
      defparam ii4231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4232 ( .DX(nn4232), .F0(dummy_35_), .F1(\cal1_u132_XORCI_8|SUM_net ), .F2(dummy_abc_2956_), .F3(dummy_abc_2957_) );
      defparam ii4232.CONFIG_DATA = 16'h8888;
      defparam ii4232.PLACE_LOCATION = "NONE";
      defparam ii4232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4233 ( .DX(nn4233), .F0(dummy_35_), .F1(\cal1_u132_XORCI_9|SUM_net ), .F2(dummy_abc_2958_), .F3(dummy_abc_2959_) );
      defparam ii4233.CONFIG_DATA = 16'h8888;
      defparam ii4233.PLACE_LOCATION = "NONE";
      defparam ii4233.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4234 ( .DX(nn4234), .F0(en), .F1(iVsyn), .F2(\coefcal1_inEn__reg|Q_net ), .F3(\coefcal1_work__reg|Q_net ) );
      defparam ii4234.CONFIG_DATA = 16'hF8F0;
      defparam ii4234.PLACE_LOCATION = "NONE";
      defparam ii4234.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4235 ( .DX(nn4235), .F0(\a_mac_out[0]_coefcal1_u64_mac_0_ ), .F1(\a_mac_out[18]_coefcal1_u64_mac ), .F2(dummy_abc_2960_), .F3(dummy_abc_2961_) );
      defparam ii4235.CONFIG_DATA = 16'h6666;
      defparam ii4235.PLACE_LOCATION = "NONE";
      defparam ii4235.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4236 ( .DX(nn4236), .F0(\a_mac_out[0]_coefcal1_u64_mac_0_ ), .F1(\a_mac_out[18]_coefcal1_u64_mac ), .F2(dummy_abc_2962_), .F3(dummy_abc_2963_) );
      defparam ii4236.CONFIG_DATA = 16'h6666;
      defparam ii4236.PLACE_LOCATION = "NONE";
      defparam ii4236.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4237 ( .DX(nn4237), .F0(\a_mac_out[19]_coefcal1_u64_mac ), .F1(\a_mac_out[1]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_2964_), .F3(dummy_abc_2965_) );
      defparam ii4237.CONFIG_DATA = 16'h6666;
      defparam ii4237.PLACE_LOCATION = "NONE";
      defparam ii4237.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4238 ( .DX(nn4238), .F0(\a_mac_out[20]_coefcal1_u64_mac ), .F1(\a_mac_out[2]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_2966_), .F3(dummy_abc_2967_) );
      defparam ii4238.CONFIG_DATA = 16'h6666;
      defparam ii4238.PLACE_LOCATION = "NONE";
      defparam ii4238.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4239 ( .DX(nn4239), .F0(\a_mac_out[21]_coefcal1_u64_mac ), .F1(\a_mac_out[3]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_2968_), .F3(dummy_abc_2969_) );
      defparam ii4239.CONFIG_DATA = 16'h6666;
      defparam ii4239.PLACE_LOCATION = "NONE";
      defparam ii4239.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4240 ( .DX(nn4240), .F0(\a_mac_out[22]_coefcal1_u64_mac ), .F1(\a_mac_out[4]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_2970_), .F3(dummy_abc_2971_) );
      defparam ii4240.CONFIG_DATA = 16'h6666;
      defparam ii4240.PLACE_LOCATION = "NONE";
      defparam ii4240.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4241 ( .DX(nn4241), .F0(\a_mac_out[23]_coefcal1_u64_mac ), .F1(\a_mac_out[5]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_2972_), .F3(dummy_abc_2973_) );
      defparam ii4241.CONFIG_DATA = 16'h6666;
      defparam ii4241.PLACE_LOCATION = "NONE";
      defparam ii4241.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4242 ( .DX(nn4242), .F0(\a_mac_out[6]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[0]_coefcal1_u64_mac ), .F2(dummy_abc_2974_), .F3(dummy_abc_2975_) );
      defparam ii4242.CONFIG_DATA = 16'h6666;
      defparam ii4242.PLACE_LOCATION = "NONE";
      defparam ii4242.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4243 ( .DX(nn4243), .F0(\a_mac_out[7]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[1]_coefcal1_u64_mac ), .F2(dummy_abc_2976_), .F3(dummy_abc_2977_) );
      defparam ii4243.CONFIG_DATA = 16'h6666;
      defparam ii4243.PLACE_LOCATION = "NONE";
      defparam ii4243.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4244 ( .DX(nn4244), .F0(\a_mac_out[8]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[2]_coefcal1_u64_mac ), .F2(dummy_abc_2978_), .F3(dummy_abc_2979_) );
      defparam ii4244.CONFIG_DATA = 16'h6666;
      defparam ii4244.PLACE_LOCATION = "NONE";
      defparam ii4244.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4245 ( .DX(nn4245), .F0(\a_mac_out[9]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[3]_coefcal1_u64_mac ), .F2(dummy_abc_2980_), .F3(dummy_abc_2981_) );
      defparam ii4245.CONFIG_DATA = 16'h6666;
      defparam ii4245.PLACE_LOCATION = "NONE";
      defparam ii4245.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4246 ( .DX(nn4246), .F0(\a_mac_out[10]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[4]_coefcal1_u64_mac ), .F2(dummy_abc_2982_), .F3(dummy_abc_2983_) );
      defparam ii4246.CONFIG_DATA = 16'h6666;
      defparam ii4246.PLACE_LOCATION = "NONE";
      defparam ii4246.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4247 ( .DX(nn4247), .F0(\a_mac_out[11]_coefcal1_u64_mac_0_ ), .F1(dummy_abc_2984_), .F2(dummy_abc_2985_), .F3(dummy_abc_2986_) );
      defparam ii4247.CONFIG_DATA = 16'hAAAA;
      defparam ii4247.PLACE_LOCATION = "NONE";
      defparam ii4247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4248 ( .DX(nn4248), .F0(\a_mac_out[12]_coefcal1_u64_mac_0_ ), .F1(dummy_abc_2987_), .F2(dummy_abc_2988_), .F3(dummy_abc_2989_) );
      defparam ii4248.CONFIG_DATA = 16'hAAAA;
      defparam ii4248.PLACE_LOCATION = "NONE";
      defparam ii4248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4249 ( .DX(nn4249), .F0(dummy_abc_2990_), .F1(dummy_abc_2991_), .F2(dummy_abc_2992_), .F3(dummy_abc_2993_) );
      defparam ii4249.CONFIG_DATA = 16'h0000;
      defparam ii4249.PLACE_LOCATION = "NONE";
      defparam ii4249.PCK_LOCATION = "NONE";
    scaler_ipc_adder_14 carry_14 ( 
        .CA( {a_acc_en_cal1_u134_mac, \a_mac_out[12]_coefcal1_u64_mac_0_ , 
              \a_mac_out[11]_coefcal1_u64_mac_0_ , \a_mac_out[10]_coefcal1_u64_mac_0_ , 
              \a_mac_out[9]_coefcal1_u64_mac_0_ , \a_mac_out[8]_coefcal1_u64_mac_0_ , 
              \a_mac_out[7]_coefcal1_u64_mac_0_ , \a_mac_out[6]_coefcal1_u64_mac_0_ , 
              \a_mac_out[5]_coefcal1_u64_mac_0_ , \a_mac_out[4]_coefcal1_u64_mac_0_ , 
              \a_mac_out[3]_coefcal1_u64_mac_0_ , \a_mac_out[2]_coefcal1_u64_mac_0_ , 
              \a_mac_out[1]_coefcal1_u64_mac_0_ , \a_mac_out[0]_coefcal1_u64_mac_0_ } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_136_ ), 
        .DX( {nn4249, nn4248, nn4247, nn4246, nn4245, nn4244, nn4243, nn4242, 
              nn4241, nn4240, nn4239, nn4238, nn4237, nn4236} ), 
        .SUM( {dummy_137_, \coefcal1_u64_XORCI_12|SUM_net , 
              \coefcal1_u64_XORCI_11|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , 
              \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u64_XORCI_8|SUM_net , 
              \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_6|SUM_net , 
              \coefcal1_u64_XORCI_5|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , 
              \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_2|SUM_net , 
              \coefcal1_u64_XORCI_1|SUM_net , \coefcal1_u64_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4266 ( .DX(nn4266), .F0(\a_mac_out[0]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[0]|Q_net ), .F2(dummy_abc_2994_), .F3(dummy_abc_2995_) );
      defparam ii4266.CONFIG_DATA = 16'h9999;
      defparam ii4266.PLACE_LOCATION = "NONE";
      defparam ii4266.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4267 ( .DX(nn4267), .F0(\a_mac_out[1]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[1]|Q_net ), .F2(dummy_abc_2996_), .F3(dummy_abc_2997_) );
      defparam ii4267.CONFIG_DATA = 16'h9999;
      defparam ii4267.PLACE_LOCATION = "NONE";
      defparam ii4267.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4268 ( .DX(nn4268), .F0(\a_mac_out[2]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[2]|Q_net ), .F2(dummy_abc_2998_), .F3(dummy_abc_2999_) );
      defparam ii4268.CONFIG_DATA = 16'h9999;
      defparam ii4268.PLACE_LOCATION = "NONE";
      defparam ii4268.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4269 ( .DX(nn4269), .F0(\a_mac_out[3]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[3]|Q_net ), .F2(dummy_abc_3000_), .F3(dummy_abc_3001_) );
      defparam ii4269.CONFIG_DATA = 16'h9999;
      defparam ii4269.PLACE_LOCATION = "NONE";
      defparam ii4269.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4270 ( .DX(nn4270), .F0(\a_mac_out[4]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[4]|Q_net ), .F2(dummy_abc_3002_), .F3(dummy_abc_3003_) );
      defparam ii4270.CONFIG_DATA = 16'h9999;
      defparam ii4270.PLACE_LOCATION = "NONE";
      defparam ii4270.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4271 ( .DX(nn4271), .F0(\a_mac_out[5]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[5]|Q_net ), .F2(dummy_abc_3004_), .F3(dummy_abc_3005_) );
      defparam ii4271.CONFIG_DATA = 16'h9999;
      defparam ii4271.PLACE_LOCATION = "NONE";
      defparam ii4271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4272 ( .DX(nn4272), .F0(\a_mac_out[6]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[6]|Q_net ), .F2(dummy_abc_3006_), .F3(dummy_abc_3007_) );
      defparam ii4272.CONFIG_DATA = 16'h9999;
      defparam ii4272.PLACE_LOCATION = "NONE";
      defparam ii4272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4273 ( .DX(nn4273), .F0(\a_mac_out[7]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[7]|Q_net ), .F2(dummy_abc_3008_), .F3(dummy_abc_3009_) );
      defparam ii4273.CONFIG_DATA = 16'h9999;
      defparam ii4273.PLACE_LOCATION = "NONE";
      defparam ii4273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4274 ( .DX(nn4274), .F0(\a_mac_out[8]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[8]|Q_net ), .F2(dummy_abc_3010_), .F3(dummy_abc_3011_) );
      defparam ii4274.CONFIG_DATA = 16'h9999;
      defparam ii4274.PLACE_LOCATION = "NONE";
      defparam ii4274.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4275 ( .DX(nn4275), .F0(\a_mac_out[9]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[9]|Q_net ), .F2(dummy_abc_3012_), .F3(dummy_abc_3013_) );
      defparam ii4275.CONFIG_DATA = 16'h9999;
      defparam ii4275.PLACE_LOCATION = "NONE";
      defparam ii4275.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4276 ( .DX(nn4276), .F0(\a_mac_out[10]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[10]|Q_net ), .F2(dummy_abc_3014_), .F3(dummy_abc_3015_) );
      defparam ii4276.CONFIG_DATA = 16'h9999;
      defparam ii4276.PLACE_LOCATION = "NONE";
      defparam ii4276.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4277 ( .DX(nn4277), .F0(\a_mac_out[11]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[11]|Q_net ), .F2(dummy_abc_3016_), .F3(dummy_abc_3017_) );
      defparam ii4277.CONFIG_DATA = 16'h9999;
      defparam ii4277.PLACE_LOCATION = "NONE";
      defparam ii4277.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4278 ( .DX(nn4278), .F0(\a_mac_out[12]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[12]|Q_net ), .F2(dummy_abc_3018_), .F3(dummy_abc_3019_) );
      defparam ii4278.CONFIG_DATA = 16'h9999;
      defparam ii4278.PLACE_LOCATION = "NONE";
      defparam ii4278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4279 ( .DX(nn4279), .F0(\a_mac_out[13]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[13]|Q_net ), .F2(dummy_abc_3020_), .F3(dummy_abc_3021_) );
      defparam ii4279.CONFIG_DATA = 16'h9999;
      defparam ii4279.PLACE_LOCATION = "NONE";
      defparam ii4279.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4280 ( .DX(nn4280), .F0(\a_mac_out[14]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[14]|Q_net ), .F2(dummy_abc_3022_), .F3(dummy_abc_3023_) );
      defparam ii4280.CONFIG_DATA = 16'h9999;
      defparam ii4280.PLACE_LOCATION = "NONE";
      defparam ii4280.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4281 ( .DX(nn4281), .F0(\a_mac_out[15]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[15]|Q_net ), .F2(dummy_abc_3024_), .F3(dummy_abc_3025_) );
      defparam ii4281.CONFIG_DATA = 16'h9999;
      defparam ii4281.PLACE_LOCATION = "NONE";
      defparam ii4281.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4282 ( .DX(nn4282), .F0(\a_mac_out[16]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[16]|Q_net ), .F2(dummy_abc_3026_), .F3(dummy_abc_3027_) );
      defparam ii4282.CONFIG_DATA = 16'h9999;
      defparam ii4282.PLACE_LOCATION = "NONE";
      defparam ii4282.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4283 ( .DX(nn4283), .F0(\a_mac_out[17]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[17]|Q_net ), .F2(dummy_abc_3028_), .F3(dummy_abc_3029_) );
      defparam ii4283.CONFIG_DATA = 16'h9999;
      defparam ii4283.PLACE_LOCATION = "NONE";
      defparam ii4283.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4284 ( .DX(nn4284), .F0(\coefcal1_working__reg[18]|Q_net ), .F1(nn4235), .F2(dummy_abc_3030_), .F3(dummy_abc_3031_) );
      defparam ii4284.CONFIG_DATA = 16'h9999;
      defparam ii4284.PLACE_LOCATION = "NONE";
      defparam ii4284.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4285 ( .DX(nn4285), .F0(\coefcal1_working__reg[19]|Q_net ), .F1(\coefcal1_u64_XORCI_1|SUM_net ), .F2(dummy_abc_3032_), .F3(dummy_abc_3033_) );
      defparam ii4285.CONFIG_DATA = 16'h9999;
      defparam ii4285.PLACE_LOCATION = "NONE";
      defparam ii4285.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4286 ( .DX(nn4286), .F0(\coefcal1_working__reg[20]|Q_net ), .F1(\coefcal1_u64_XORCI_2|SUM_net ), .F2(dummy_abc_3034_), .F3(dummy_abc_3035_) );
      defparam ii4286.CONFIG_DATA = 16'h9999;
      defparam ii4286.PLACE_LOCATION = "NONE";
      defparam ii4286.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4287 ( .DX(nn4287), .F0(\coefcal1_working__reg[21]|Q_net ), .F1(\coefcal1_u64_XORCI_3|SUM_net ), .F2(dummy_abc_3036_), .F3(dummy_abc_3037_) );
      defparam ii4287.CONFIG_DATA = 16'h9999;
      defparam ii4287.PLACE_LOCATION = "NONE";
      defparam ii4287.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4288 ( .DX(nn4288), .F0(\coefcal1_working__reg[22]|Q_net ), .F1(\coefcal1_u64_XORCI_4|SUM_net ), .F2(dummy_abc_3038_), .F3(dummy_abc_3039_) );
      defparam ii4288.CONFIG_DATA = 16'h9999;
      defparam ii4288.PLACE_LOCATION = "NONE";
      defparam ii4288.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4289 ( .DX(nn4289), .F0(\coefcal1_working__reg[23]|Q_net ), .F1(\coefcal1_u64_XORCI_5|SUM_net ), .F2(dummy_abc_3040_), .F3(dummy_abc_3041_) );
      defparam ii4289.CONFIG_DATA = 16'h9999;
      defparam ii4289.PLACE_LOCATION = "NONE";
      defparam ii4289.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4290 ( .DX(nn4290), .F0(\coefcal1_working__reg[24]|Q_net ), .F1(\coefcal1_u64_XORCI_6|SUM_net ), .F2(dummy_abc_3042_), .F3(dummy_abc_3043_) );
      defparam ii4290.CONFIG_DATA = 16'h9999;
      defparam ii4290.PLACE_LOCATION = "NONE";
      defparam ii4290.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4291 ( .DX(nn4291), .F0(\coefcal1_working__reg[25]|Q_net ), .F1(\coefcal1_u64_XORCI_7|SUM_net ), .F2(dummy_abc_3044_), .F3(dummy_abc_3045_) );
      defparam ii4291.CONFIG_DATA = 16'h9999;
      defparam ii4291.PLACE_LOCATION = "NONE";
      defparam ii4291.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4292 ( .DX(nn4292), .F0(\coefcal1_working__reg[26]|Q_net ), .F1(\coefcal1_u64_XORCI_8|SUM_net ), .F2(dummy_abc_3046_), .F3(dummy_abc_3047_) );
      defparam ii4292.CONFIG_DATA = 16'h9999;
      defparam ii4292.PLACE_LOCATION = "NONE";
      defparam ii4292.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4293 ( .DX(nn4293), .F0(\coefcal1_working__reg[27]|Q_net ), .F1(\coefcal1_u64_XORCI_9|SUM_net ), .F2(dummy_abc_3048_), .F3(dummy_abc_3049_) );
      defparam ii4293.CONFIG_DATA = 16'h9999;
      defparam ii4293.PLACE_LOCATION = "NONE";
      defparam ii4293.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4294 ( .DX(nn4294), .F0(\coefcal1_working__reg[28]|Q_net ), .F1(\coefcal1_u64_XORCI_10|SUM_net ), .F2(dummy_abc_3050_), .F3(dummy_abc_3051_) );
      defparam ii4294.CONFIG_DATA = 16'h9999;
      defparam ii4294.PLACE_LOCATION = "NONE";
      defparam ii4294.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4295 ( .DX(nn4295), .F0(\coefcal1_working__reg[29]|Q_net ), .F1(\coefcal1_u64_XORCI_11|SUM_net ), .F2(dummy_abc_3052_), .F3(dummy_abc_3053_) );
      defparam ii4295.CONFIG_DATA = 16'h9999;
      defparam ii4295.PLACE_LOCATION = "NONE";
      defparam ii4295.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4296 ( .DX(nn4296), .F0(\coefcal1_working__reg[30]|Q_net ), .F1(\coefcal1_u64_XORCI_12|SUM_net ), .F2(dummy_abc_3054_), .F3(dummy_abc_3055_) );
      defparam ii4296.CONFIG_DATA = 16'h9999;
      defparam ii4296.PLACE_LOCATION = "NONE";
      defparam ii4296.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4297 ( .DX(nn4297), .F0(\coefcal1_working__reg[31]|Q_net ), .F1(dummy_abc_3056_), .F2(dummy_abc_3057_), .F3(dummy_abc_3058_) );
      defparam ii4297.CONFIG_DATA = 16'h5555;
      defparam ii4297.PLACE_LOCATION = "NONE";
      defparam ii4297.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4298 ( .DX(nn4298), .F0(\coefcal1_working__reg[32]|Q_net ), .F1(dummy_abc_3059_), .F2(dummy_abc_3060_), .F3(dummy_abc_3061_) );
      defparam ii4298.CONFIG_DATA = 16'h5555;
      defparam ii4298.PLACE_LOCATION = "NONE";
      defparam ii4298.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4299 ( .DX(nn4299), .F0(dummy_abc_3062_), .F1(dummy_abc_3063_), .F2(dummy_abc_3064_), .F3(dummy_abc_3065_) );
      defparam ii4299.CONFIG_DATA = 16'hFFFF;
      defparam ii4299.PLACE_LOCATION = "NONE";
      defparam ii4299.PCK_LOCATION = "NONE";
    scaler_ipc_adder_34 carry_34 ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, \coefcal1_u64_XORCI_12|SUM_net , 
              \coefcal1_u64_XORCI_11|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , 
              \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u64_XORCI_8|SUM_net , 
              \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_6|SUM_net , 
              \coefcal1_u64_XORCI_5|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , 
              \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_2|SUM_net , 
              \coefcal1_u64_XORCI_1|SUM_net , nn4235, \a_mac_out[17]_coefcal1_u64_mac , 
              \a_mac_out[16]_coefcal1_u64_mac , \a_mac_out[15]_coefcal1_u64_mac , 
              \a_mac_out[14]_coefcal1_u64_mac , \a_mac_out[13]_coefcal1_u64_mac , 
              \a_mac_out[12]_coefcal1_u64_mac , \a_mac_out[11]_coefcal1_u64_mac , 
              \a_mac_out[10]_coefcal1_u64_mac , \a_mac_out[9]_coefcal1_u64_mac , 
              \a_mac_out[8]_coefcal1_u64_mac , \a_mac_out[7]_coefcal1_u64_mac , 
              \a_mac_out[6]_coefcal1_u64_mac , \a_mac_out[5]_coefcal1_u64_mac , 
              \a_mac_out[4]_coefcal1_u64_mac , \a_mac_out[3]_coefcal1_u64_mac , 
              \a_mac_out[2]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u64_mac , 
              \a_mac_out[0]_coefcal1_u64_mac } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_849_ ), 
        .DX( {nn4299, nn4298, nn4297, nn4296, nn4295, nn4294, nn4293, nn4292, 
              nn4291, nn4290, nn4289, nn4288, nn4287, nn4286, nn4285, nn4284, 
              nn4283, nn4282, nn4281, nn4280, nn4279, nn4278, nn4277, nn4276, 
              nn4275, nn4274, nn4273, nn4272, nn4271, nn4270, nn4269, nn4268, 
              nn4267, nn4266} ), 
        .SUM( {\coefcal1_u8_XORCI_33|SUM_net , dummy_850_, dummy_851_, dummy_852_, 
              dummy_853_, dummy_854_, dummy_855_, dummy_856_, dummy_857_, dummy_858_, 
              dummy_859_, dummy_860_, dummy_861_, dummy_862_, dummy_863_, dummy_864_, 
              dummy_865_, dummy_866_, dummy_867_, dummy_868_, dummy_869_, dummy_870_, 
              dummy_871_, dummy_872_, dummy_873_, dummy_874_, dummy_875_, dummy_876_, 
              dummy_877_, dummy_878_, dummy_879_, dummy_880_, dummy_881_, dummy_882_} )
      );
    CS_LUT4_PRIM ii4336 ( .DX(nn4336), .F0(dummy_849_), .F1(dummy_abc_3066_), .F2(dummy_abc_3067_), .F3(dummy_abc_3068_) );
      defparam ii4336.CONFIG_DATA = 16'h5555;
      defparam ii4336.PLACE_LOCATION = "NONE";
      defparam ii4336.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4337 ( .DX(nn4337), .F0(nn0812), .F1(dummy_abc_3069_), .F2(dummy_abc_3070_), .F3(dummy_abc_3071_) );
      defparam ii4337.CONFIG_DATA = 16'h5555;
      defparam ii4337.PLACE_LOCATION = "NONE";
      defparam ii4337.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4338 ( .DX(nn4338), .F0(\u2_XORCI_1|SUM_net ), .F1(dummy_abc_3072_), .F2(dummy_abc_3073_), .F3(dummy_abc_3074_) );
      defparam ii4338.CONFIG_DATA = 16'hAAAA;
      defparam ii4338.PLACE_LOCATION = "NONE";
      defparam ii4338.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4339 ( .DX(nn4339), .F0(\u2_XORCI_2|SUM_net ), .F1(dummy_abc_3075_), .F2(dummy_abc_3076_), .F3(dummy_abc_3077_) );
      defparam ii4339.CONFIG_DATA = 16'hAAAA;
      defparam ii4339.PLACE_LOCATION = "NONE";
      defparam ii4339.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4340 ( .DX(nn4340), .F0(\u2_XORCI_3|SUM_net ), .F1(dummy_abc_3078_), .F2(dummy_abc_3079_), .F3(dummy_abc_3080_) );
      defparam ii4340.CONFIG_DATA = 16'hAAAA;
      defparam ii4340.PLACE_LOCATION = "NONE";
      defparam ii4340.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4341 ( .DX(nn4341), .F0(\u2_XORCI_4|SUM_net ), .F1(dummy_abc_3081_), .F2(dummy_abc_3082_), .F3(dummy_abc_3083_) );
      defparam ii4341.CONFIG_DATA = 16'hAAAA;
      defparam ii4341.PLACE_LOCATION = "NONE";
      defparam ii4341.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4342 ( .DX(nn4342), .F0(\u2_XORCI_5|SUM_net ), .F1(dummy_abc_3084_), .F2(dummy_abc_3085_), .F3(dummy_abc_3086_) );
      defparam ii4342.CONFIG_DATA = 16'hAAAA;
      defparam ii4342.PLACE_LOCATION = "NONE";
      defparam ii4342.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4343 ( .DX(nn4343), .F0(\u2_XORCI_6|SUM_net ), .F1(dummy_abc_3087_), .F2(dummy_abc_3088_), .F3(dummy_abc_3089_) );
      defparam ii4343.CONFIG_DATA = 16'hAAAA;
      defparam ii4343.PLACE_LOCATION = "NONE";
      defparam ii4343.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4344 ( .DX(nn4344), .F0(\u2_XORCI_7|SUM_net ), .F1(dummy_abc_3090_), .F2(dummy_abc_3091_), .F3(dummy_abc_3092_) );
      defparam ii4344.CONFIG_DATA = 16'hAAAA;
      defparam ii4344.PLACE_LOCATION = "NONE";
      defparam ii4344.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4345 ( .DX(nn4345), .F0(\u2_XORCI_8|SUM_net ), .F1(dummy_abc_3093_), .F2(dummy_abc_3094_), .F3(dummy_abc_3095_) );
      defparam ii4345.CONFIG_DATA = 16'hAAAA;
      defparam ii4345.PLACE_LOCATION = "NONE";
      defparam ii4345.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4346 ( .DX(nn4346), .F0(\u2_XORCI_9|SUM_net ), .F1(dummy_abc_3096_), .F2(dummy_abc_3097_), .F3(dummy_abc_3098_) );
      defparam ii4346.CONFIG_DATA = 16'hAAAA;
      defparam ii4346.PLACE_LOCATION = "NONE";
      defparam ii4346.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4347 ( .DX(nn4347), .F0(\u2_XORCI_10|SUM_net ), .F1(dummy_abc_3099_), .F2(dummy_abc_3100_), .F3(dummy_abc_3101_) );
      defparam ii4347.CONFIG_DATA = 16'hAAAA;
      defparam ii4347.PLACE_LOCATION = "NONE";
      defparam ii4347.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_72_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_dinxy_cen_cal1_u134_mac} ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_16_ ), 
        .DX( {nn4347, nn4346, nn4345, nn4344, nn4343, nn4342, nn4341, nn4340, 
              nn4339, nn4338, nn4337} ), 
        .SUM( {\coefcal1_u59_XORCI_10|SUM_net , \coefcal1_u59_XORCI_9|SUM_net , 
              \coefcal1_u59_XORCI_8|SUM_net , \coefcal1_u59_XORCI_7|SUM_net , 
              \coefcal1_u59_XORCI_6|SUM_net , \coefcal1_u59_XORCI_5|SUM_net , 
              \coefcal1_u59_XORCI_4|SUM_net , \coefcal1_u59_XORCI_3|SUM_net , 
              \coefcal1_u59_XORCI_2|SUM_net , \coefcal1_u59_XORCI_1|SUM_net , 
              \coefcal1_u59_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4361 ( .DX(nn4361), .F0(nn0812), .F1(dummy_abc_3102_), .F2(dummy_abc_3103_), .F3(dummy_abc_3104_) );
      defparam ii4361.CONFIG_DATA = 16'h5555;
      defparam ii4361.PLACE_LOCATION = "NONE";
      defparam ii4361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4362 ( .DX(nn4362), .F0(\u3_XORCI_1|SUM_net ), .F1(dummy_abc_3105_), .F2(dummy_abc_3106_), .F3(dummy_abc_3107_) );
      defparam ii4362.CONFIG_DATA = 16'h5555;
      defparam ii4362.PLACE_LOCATION = "NONE";
      defparam ii4362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4363 ( .DX(nn4363), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3108_), .F3(dummy_abc_3109_) );
      defparam ii4363.CONFIG_DATA = 16'h9999;
      defparam ii4363.PLACE_LOCATION = "NONE";
      defparam ii4363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4364 ( .DX(nn4364), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3110_), .F3(dummy_abc_3111_) );
      defparam ii4364.CONFIG_DATA = 16'h9999;
      defparam ii4364.PLACE_LOCATION = "NONE";
      defparam ii4364.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4365 ( .DX(nn4365), .F0(yBgn[1]), .F1(yEnd[1]), .F2(dummy_abc_3112_), .F3(dummy_abc_3113_) );
      defparam ii4365.CONFIG_DATA = 16'h9999;
      defparam ii4365.PLACE_LOCATION = "NONE";
      defparam ii4365.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4366 ( .DX(nn4366), .F0(yBgn[2]), .F1(yEnd[2]), .F2(dummy_abc_3114_), .F3(dummy_abc_3115_) );
      defparam ii4366.CONFIG_DATA = 16'h9999;
      defparam ii4366.PLACE_LOCATION = "NONE";
      defparam ii4366.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4367 ( .DX(nn4367), .F0(yBgn[3]), .F1(yEnd[3]), .F2(dummy_abc_3116_), .F3(dummy_abc_3117_) );
      defparam ii4367.CONFIG_DATA = 16'h9999;
      defparam ii4367.PLACE_LOCATION = "NONE";
      defparam ii4367.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4368 ( .DX(nn4368), .F0(yBgn[4]), .F1(yEnd[4]), .F2(dummy_abc_3118_), .F3(dummy_abc_3119_) );
      defparam ii4368.CONFIG_DATA = 16'h9999;
      defparam ii4368.PLACE_LOCATION = "NONE";
      defparam ii4368.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4369 ( .DX(nn4369), .F0(yBgn[5]), .F1(yEnd[5]), .F2(dummy_abc_3120_), .F3(dummy_abc_3121_) );
      defparam ii4369.CONFIG_DATA = 16'h9999;
      defparam ii4369.PLACE_LOCATION = "NONE";
      defparam ii4369.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4370 ( .DX(nn4370), .F0(yBgn[6]), .F1(yEnd[6]), .F2(dummy_abc_3122_), .F3(dummy_abc_3123_) );
      defparam ii4370.CONFIG_DATA = 16'h9999;
      defparam ii4370.PLACE_LOCATION = "NONE";
      defparam ii4370.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4371 ( .DX(nn4371), .F0(yBgn[7]), .F1(yEnd[7]), .F2(dummy_abc_3124_), .F3(dummy_abc_3125_) );
      defparam ii4371.CONFIG_DATA = 16'h9999;
      defparam ii4371.PLACE_LOCATION = "NONE";
      defparam ii4371.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4372 ( .DX(nn4372), .F0(yBgn[8]), .F1(yEnd[8]), .F2(dummy_abc_3126_), .F3(dummy_abc_3127_) );
      defparam ii4372.CONFIG_DATA = 16'h9999;
      defparam ii4372.PLACE_LOCATION = "NONE";
      defparam ii4372.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4373 ( .DX(nn4373), .F0(yBgn[9]), .F1(yEnd[9]), .F2(dummy_abc_3128_), .F3(dummy_abc_3129_) );
      defparam ii4373.CONFIG_DATA = 16'h9999;
      defparam ii4373.PLACE_LOCATION = "NONE";
      defparam ii4373.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4374 ( .DX(nn4374), .F0(yBgn[10]), .F1(yEnd[10]), .F2(dummy_abc_3130_), .F3(dummy_abc_3131_) );
      defparam ii4374.CONFIG_DATA = 16'h9999;
      defparam ii4374.PLACE_LOCATION = "NONE";
      defparam ii4374.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4375 ( .DX(nn4375), .F0(dummy_abc_3132_), .F1(dummy_abc_3133_), .F2(dummy_abc_3134_), .F3(dummy_abc_3135_) );
      defparam ii4375.CONFIG_DATA = 16'hFFFF;
      defparam ii4375.PLACE_LOCATION = "NONE";
      defparam ii4375.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_76_ ( 
        .CA( {a_acc_en_cal1_u134_mac, yEnd[10], yEnd[9], yEnd[8], yEnd[7], 
              yEnd[6], yEnd[5], yEnd[4], yEnd[3], yEnd[2], yEnd[1], yEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_49_ ), 
        .DX( {nn4375, nn4374, nn4373, nn4372, nn4371, nn4370, nn4369, nn4368, 
              nn4367, nn4366, nn4365, nn4364} ), 
        .SUM( {dummy_50_, \coefcal1_u7_XORCI_10|SUM_net , 
              \coefcal1_u7_XORCI_9|SUM_net , \coefcal1_u7_XORCI_8|SUM_net , 
              \coefcal1_u7_XORCI_7|SUM_net , \coefcal1_u7_XORCI_6|SUM_net , 
              \coefcal1_u7_XORCI_5|SUM_net , \coefcal1_u7_XORCI_4|SUM_net , 
              \coefcal1_u7_XORCI_3|SUM_net , \coefcal1_u7_XORCI_2|SUM_net , 
              \coefcal1_u7_XORCI_1|SUM_net , \coefcal1_u7_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4390 ( .DX(nn4390), .F0(\coefcal1_u7_XORCI_1|SUM_net ), .F1(dummy_abc_3136_), .F2(dummy_abc_3137_), .F3(dummy_abc_3138_) );
      defparam ii4390.CONFIG_DATA = 16'hAAAA;
      defparam ii4390.PLACE_LOCATION = "NONE";
      defparam ii4390.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4391 ( .DX(nn4391), .F0(\coefcal1_u7_XORCI_2|SUM_net ), .F1(dummy_abc_3139_), .F2(dummy_abc_3140_), .F3(dummy_abc_3141_) );
      defparam ii4391.CONFIG_DATA = 16'hAAAA;
      defparam ii4391.PLACE_LOCATION = "NONE";
      defparam ii4391.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4392 ( .DX(nn4392), .F0(\coefcal1_u7_XORCI_3|SUM_net ), .F1(dummy_abc_3142_), .F2(dummy_abc_3143_), .F3(dummy_abc_3144_) );
      defparam ii4392.CONFIG_DATA = 16'hAAAA;
      defparam ii4392.PLACE_LOCATION = "NONE";
      defparam ii4392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4393 ( .DX(nn4393), .F0(\coefcal1_u7_XORCI_4|SUM_net ), .F1(dummy_abc_3145_), .F2(dummy_abc_3146_), .F3(dummy_abc_3147_) );
      defparam ii4393.CONFIG_DATA = 16'hAAAA;
      defparam ii4393.PLACE_LOCATION = "NONE";
      defparam ii4393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4394 ( .DX(nn4394), .F0(\coefcal1_u7_XORCI_5|SUM_net ), .F1(dummy_abc_3148_), .F2(dummy_abc_3149_), .F3(dummy_abc_3150_) );
      defparam ii4394.CONFIG_DATA = 16'hAAAA;
      defparam ii4394.PLACE_LOCATION = "NONE";
      defparam ii4394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4395 ( .DX(nn4395), .F0(\coefcal1_u7_XORCI_6|SUM_net ), .F1(dummy_abc_3151_), .F2(dummy_abc_3152_), .F3(dummy_abc_3153_) );
      defparam ii4395.CONFIG_DATA = 16'hAAAA;
      defparam ii4395.PLACE_LOCATION = "NONE";
      defparam ii4395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4396 ( .DX(nn4396), .F0(\coefcal1_u7_XORCI_7|SUM_net ), .F1(dummy_abc_3154_), .F2(dummy_abc_3155_), .F3(dummy_abc_3156_) );
      defparam ii4396.CONFIG_DATA = 16'hAAAA;
      defparam ii4396.PLACE_LOCATION = "NONE";
      defparam ii4396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4397 ( .DX(nn4397), .F0(\coefcal1_u7_XORCI_8|SUM_net ), .F1(dummy_abc_3157_), .F2(dummy_abc_3158_), .F3(dummy_abc_3159_) );
      defparam ii4397.CONFIG_DATA = 16'hAAAA;
      defparam ii4397.PLACE_LOCATION = "NONE";
      defparam ii4397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4398 ( .DX(nn4398), .F0(\coefcal1_u7_XORCI_9|SUM_net ), .F1(dummy_abc_3160_), .F2(dummy_abc_3161_), .F3(dummy_abc_3162_) );
      defparam ii4398.CONFIG_DATA = 16'hAAAA;
      defparam ii4398.PLACE_LOCATION = "NONE";
      defparam ii4398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4399 ( .DX(nn4399), .F0(\coefcal1_u7_XORCI_10|SUM_net ), .F1(dummy_abc_3163_), .F2(dummy_abc_3164_), .F3(dummy_abc_3165_) );
      defparam ii4399.CONFIG_DATA = 16'hAAAA;
      defparam ii4399.PLACE_LOCATION = "NONE";
      defparam ii4399.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_73_ ( 
        .CA( {a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, 
              a_acc_en_cal1_u134_mac, a_acc_en_cal1_u134_mac, a_dinxy_cen_cal1_u134_mac} ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_17_ ), 
        .DX( {nn4399, nn4398, nn4397, nn4396, nn4395, nn4394, nn4393, nn4392, 
              nn4391, nn4390, nn4363} ), 
        .SUM( {\coefcal1_u60_XORCI_10|SUM_net , \coefcal1_u60_XORCI_9|SUM_net , 
              \coefcal1_u60_XORCI_8|SUM_net , \coefcal1_u60_XORCI_7|SUM_net , 
              \coefcal1_u60_XORCI_6|SUM_net , \coefcal1_u60_XORCI_5|SUM_net , 
              \coefcal1_u60_XORCI_4|SUM_net , \coefcal1_u60_XORCI_3|SUM_net , 
              \coefcal1_u60_XORCI_2|SUM_net , \coefcal1_u60_XORCI_1|SUM_net , 
              \coefcal1_u60_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4413 ( .DX(nn4413), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3166_), .F3(dummy_abc_3167_) );
      defparam ii4413.CONFIG_DATA = 16'h9999;
      defparam ii4413.PLACE_LOCATION = "NONE";
      defparam ii4413.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4414 ( .DX(nn4414), .F0(dIn[0]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3168_) );
      defparam ii4414.CONFIG_DATA = 16'h0202;
      defparam ii4414.PLACE_LOCATION = "NONE";
      defparam ii4414.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4415 ( .DX(nn4415), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(\inputctrl1_yAddress__reg[1]|Q_net ), .F2(\inputctrl1_yCal__reg[6]|Q_net ), .F3(\inputctrl1_yCal__reg[7]|Q_net ) );
      defparam ii4415.CONFIG_DATA = 16'h8421;
      defparam ii4415.PLACE_LOCATION = "NONE";
      defparam ii4415.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4416 ( .DX(nn4416), .F0(\inputctrl1_yAddress__reg[5]|Q_net ), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(\inputctrl1_yCal__reg[11]|Q_net ), .F3(\inputctrl1_yCal__reg[14]|Q_net ) );
      defparam ii4416.CONFIG_DATA = 16'h8421;
      defparam ii4416.PLACE_LOCATION = "NONE";
      defparam ii4416.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4417 ( .DX(nn4417), .F0(\inputctrl1_yAddress__reg[3]|Q_net ), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(\inputctrl1_yCal__reg[15]|Q_net ), .F3(\inputctrl1_yCal__reg[9]|Q_net ) );
      defparam ii4417.CONFIG_DATA = 16'h8241;
      defparam ii4417.PLACE_LOCATION = "NONE";
      defparam ii4417.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4418 ( .DX(nn4418), .F0(\inputctrl1_yAddress__reg[10]|Q_net ), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(\inputctrl1_yCal__reg[13]|Q_net ), .F3(\inputctrl1_yCal__reg[16]|Q_net ) );
      defparam ii4418.CONFIG_DATA = 16'h8241;
      defparam ii4418.PLACE_LOCATION = "NONE";
      defparam ii4418.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4419 ( .DX(nn4419), .F0(\inputctrl1_yAddress__reg[2]|Q_net ), .F1(\inputctrl1_yAddress__reg[4]|Q_net ), .F2(\inputctrl1_yCal__reg[10]|Q_net ), .F3(\inputctrl1_yCal__reg[8]|Q_net ) );
      defparam ii4419.CONFIG_DATA = 16'h8241;
      defparam ii4419.PLACE_LOCATION = "NONE";
      defparam ii4419.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4420 ( .DX(nn4420), .F0(nn4416), .F1(nn4417), .F2(nn4418), .F3(nn4419) );
      defparam ii4420.CONFIG_DATA = 16'h8000;
      defparam ii4420.PLACE_LOCATION = "NONE";
      defparam ii4420.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4421 ( .DX(nn4421), .F0(\inputctrl1_yAddress__reg[6]|Q_net ), .F1(\inputctrl1_yCal__reg[12]|Q_net ), .F2(nn4415), .F3(nn4420) );
      defparam ii4421.CONFIG_DATA = 16'h9000;
      defparam ii4421.PLACE_LOCATION = "NONE";
      defparam ii4421.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4422 ( .DX(nn4422), .F0(\inputctrl1_yPreEn__reg|Q_net ), .F1(nn4421), .F2(dummy_abc_3169_), .F3(dummy_abc_3170_) );
      defparam ii4422.CONFIG_DATA = 16'h1111;
      defparam ii4422.PLACE_LOCATION = "NONE";
      defparam ii4422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4423 ( .DX(nn4423), .F0(yEnd[0]), .F1(\inputctrl1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_3171_), .F3(dummy_abc_3172_) );
      defparam ii4423.CONFIG_DATA = 16'h9999;
      defparam ii4423.PLACE_LOCATION = "NONE";
      defparam ii4423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4424 ( .DX(nn4424), .F0(yEnd[1]), .F1(\inputctrl1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_3173_), .F3(dummy_abc_3174_) );
      defparam ii4424.CONFIG_DATA = 16'h9999;
      defparam ii4424.PLACE_LOCATION = "NONE";
      defparam ii4424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4425 ( .DX(nn4425), .F0(yEnd[2]), .F1(\inputctrl1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_3175_), .F3(dummy_abc_3176_) );
      defparam ii4425.CONFIG_DATA = 16'h9999;
      defparam ii4425.PLACE_LOCATION = "NONE";
      defparam ii4425.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4426 ( .DX(nn4426), .F0(yEnd[3]), .F1(\inputctrl1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_3177_), .F3(dummy_abc_3178_) );
      defparam ii4426.CONFIG_DATA = 16'h9999;
      defparam ii4426.PLACE_LOCATION = "NONE";
      defparam ii4426.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4427 ( .DX(nn4427), .F0(yEnd[4]), .F1(\inputctrl1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_3179_), .F3(dummy_abc_3180_) );
      defparam ii4427.CONFIG_DATA = 16'h9999;
      defparam ii4427.PLACE_LOCATION = "NONE";
      defparam ii4427.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4428 ( .DX(nn4428), .F0(yEnd[5]), .F1(\inputctrl1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_3181_), .F3(dummy_abc_3182_) );
      defparam ii4428.CONFIG_DATA = 16'h9999;
      defparam ii4428.PLACE_LOCATION = "NONE";
      defparam ii4428.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4429 ( .DX(nn4429), .F0(yEnd[6]), .F1(\inputctrl1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_3183_), .F3(dummy_abc_3184_) );
      defparam ii4429.CONFIG_DATA = 16'h9999;
      defparam ii4429.PLACE_LOCATION = "NONE";
      defparam ii4429.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4430 ( .DX(nn4430), .F0(yEnd[7]), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_3185_), .F3(dummy_abc_3186_) );
      defparam ii4430.CONFIG_DATA = 16'h9999;
      defparam ii4430.PLACE_LOCATION = "NONE";
      defparam ii4430.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4431 ( .DX(nn4431), .F0(yEnd[8]), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_3187_), .F3(dummy_abc_3188_) );
      defparam ii4431.CONFIG_DATA = 16'h9999;
      defparam ii4431.PLACE_LOCATION = "NONE";
      defparam ii4431.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4432 ( .DX(nn4432), .F0(yEnd[9]), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_3189_), .F3(dummy_abc_3190_) );
      defparam ii4432.CONFIG_DATA = 16'h9999;
      defparam ii4432.PLACE_LOCATION = "NONE";
      defparam ii4432.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4433 ( .DX(nn4433), .F0(yEnd[10]), .F1(\inputctrl1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_3191_), .F3(dummy_abc_3192_) );
      defparam ii4433.CONFIG_DATA = 16'h9999;
      defparam ii4433.PLACE_LOCATION = "NONE";
      defparam ii4433.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4434 ( .DX(nn4434), .F0(dummy_abc_3193_), .F1(dummy_abc_3194_), .F2(dummy_abc_3195_), .F3(dummy_abc_3196_) );
      defparam ii4434.CONFIG_DATA = 16'hFFFF;
      defparam ii4434.PLACE_LOCATION = "NONE";
      defparam ii4434.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_85_ ( 
        .CA( {a_acc_en_cal1_u134_mac, yEnd[10], yEnd[9], yEnd[8], yEnd[7], 
              yEnd[6], yEnd[5], yEnd[4], yEnd[3], yEnd[2], yEnd[1], yEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_104_ ), 
        .DX( {nn4434, nn4433, nn4432, nn4431, nn4430, nn4429, nn4428, nn4427, 
              nn4426, nn4425, nn4424, nn4423} ), 
        .SUM( {\inputctrl1_u43_XORCI_11|SUM_net , dummy_105_, dummy_106_, 
              dummy_107_, dummy_108_, dummy_109_, dummy_110_, dummy_111_, dummy_112_, 
              dummy_113_, dummy_114_, dummy_115_} )
      );
    CS_LUT4_PRIM ii4449 ( .DX(nn4449), .F0(\inputctrl1_xAddress__reg[3]|Q_net ), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(\inputctrl1_xCal__reg[12]|Q_net ), .F3(\inputctrl1_xCal__reg[9]|Q_net ) );
      defparam ii4449.CONFIG_DATA = 16'h8241;
      defparam ii4449.PLACE_LOCATION = "NONE";
      defparam ii4449.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4450 ( .DX(nn4450), .F0(\inputctrl1_xAddress__reg[1]|Q_net ), .F1(\inputctrl1_xAddress__reg[2]|Q_net ), .F2(\inputctrl1_xCal__reg[7]|Q_net ), .F3(\inputctrl1_xCal__reg[8]|Q_net ) );
      defparam ii4450.CONFIG_DATA = 16'h8421;
      defparam ii4450.PLACE_LOCATION = "NONE";
      defparam ii4450.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4451 ( .DX(nn4451), .F0(\inputctrl1_xAddress__reg[4]|Q_net ), .F1(\inputctrl1_xAddress__reg[7]|Q_net ), .F2(\inputctrl1_xCal__reg[10]|Q_net ), .F3(\inputctrl1_xCal__reg[13]|Q_net ) );
      defparam ii4451.CONFIG_DATA = 16'h8421;
      defparam ii4451.PLACE_LOCATION = "NONE";
      defparam ii4451.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4452 ( .DX(nn4452), .F0(\inputctrl1_xAddress__reg[5]|Q_net ), .F1(\inputctrl1_xAddress__reg[8]|Q_net ), .F2(\inputctrl1_xCal__reg[11]|Q_net ), .F3(\inputctrl1_xCal__reg[14]|Q_net ) );
      defparam ii4452.CONFIG_DATA = 16'h8421;
      defparam ii4452.PLACE_LOCATION = "NONE";
      defparam ii4452.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4453 ( .DX(nn4453), .F0(nn4449), .F1(nn4450), .F2(nn4451), .F3(nn4452) );
      defparam ii4453.CONFIG_DATA = 16'h8000;
      defparam ii4453.PLACE_LOCATION = "NONE";
      defparam ii4453.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4454 ( .DX(nn4454), .F0(\inputctrl1_xAddress__reg[10]|Q_net ), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(\inputctrl1_xCal__reg[15]|Q_net ), .F3(\inputctrl1_xCal__reg[16]|Q_net ) );
      defparam ii4454.CONFIG_DATA = 16'h8241;
      defparam ii4454.PLACE_LOCATION = "NONE";
      defparam ii4454.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4455 ( .DX(nn4455), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(\inputctrl1_xCal__reg[6]|Q_net ), .F2(nn4453), .F3(nn4454) );
      defparam ii4455.CONFIG_DATA = 16'h9000;
      defparam ii4455.PLACE_LOCATION = "NONE";
      defparam ii4455.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4456 ( .DX(nn4456), .F0(xEnd[0]), .F1(\inputctrl1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_3197_), .F3(dummy_abc_3198_) );
      defparam ii4456.CONFIG_DATA = 16'h9999;
      defparam ii4456.PLACE_LOCATION = "NONE";
      defparam ii4456.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4457 ( .DX(nn4457), .F0(xEnd[1]), .F1(\inputctrl1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_3199_), .F3(dummy_abc_3200_) );
      defparam ii4457.CONFIG_DATA = 16'h9999;
      defparam ii4457.PLACE_LOCATION = "NONE";
      defparam ii4457.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4458 ( .DX(nn4458), .F0(xEnd[2]), .F1(\inputctrl1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_3201_), .F3(dummy_abc_3202_) );
      defparam ii4458.CONFIG_DATA = 16'h9999;
      defparam ii4458.PLACE_LOCATION = "NONE";
      defparam ii4458.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4459 ( .DX(nn4459), .F0(xEnd[3]), .F1(\inputctrl1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_3203_), .F3(dummy_abc_3204_) );
      defparam ii4459.CONFIG_DATA = 16'h9999;
      defparam ii4459.PLACE_LOCATION = "NONE";
      defparam ii4459.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4460 ( .DX(nn4460), .F0(xEnd[4]), .F1(\inputctrl1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_3205_), .F3(dummy_abc_3206_) );
      defparam ii4460.CONFIG_DATA = 16'h9999;
      defparam ii4460.PLACE_LOCATION = "NONE";
      defparam ii4460.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4461 ( .DX(nn4461), .F0(xEnd[5]), .F1(\inputctrl1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_3207_), .F3(dummy_abc_3208_) );
      defparam ii4461.CONFIG_DATA = 16'h9999;
      defparam ii4461.PLACE_LOCATION = "NONE";
      defparam ii4461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4462 ( .DX(nn4462), .F0(xEnd[6]), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_3209_), .F3(dummy_abc_3210_) );
      defparam ii4462.CONFIG_DATA = 16'h9999;
      defparam ii4462.PLACE_LOCATION = "NONE";
      defparam ii4462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4463 ( .DX(nn4463), .F0(xEnd[7]), .F1(\inputctrl1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_3211_), .F3(dummy_abc_3212_) );
      defparam ii4463.CONFIG_DATA = 16'h9999;
      defparam ii4463.PLACE_LOCATION = "NONE";
      defparam ii4463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4464 ( .DX(nn4464), .F0(xEnd[8]), .F1(\inputctrl1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_3213_), .F3(dummy_abc_3214_) );
      defparam ii4464.CONFIG_DATA = 16'h9999;
      defparam ii4464.PLACE_LOCATION = "NONE";
      defparam ii4464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4465 ( .DX(nn4465), .F0(xEnd[9]), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_3215_), .F3(dummy_abc_3216_) );
      defparam ii4465.CONFIG_DATA = 16'h9999;
      defparam ii4465.PLACE_LOCATION = "NONE";
      defparam ii4465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4466 ( .DX(nn4466), .F0(xEnd[10]), .F1(\inputctrl1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_3217_), .F3(dummy_abc_3218_) );
      defparam ii4466.CONFIG_DATA = 16'h9999;
      defparam ii4466.PLACE_LOCATION = "NONE";
      defparam ii4466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4467 ( .DX(nn4467), .F0(dummy_abc_3219_), .F1(dummy_abc_3220_), .F2(dummy_abc_3221_), .F3(dummy_abc_3222_) );
      defparam ii4467.CONFIG_DATA = 16'hFFFF;
      defparam ii4467.PLACE_LOCATION = "NONE";
      defparam ii4467.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_84_ ( 
        .CA( {a_acc_en_cal1_u134_mac, xEnd[10], xEnd[9], xEnd[8], xEnd[7], 
              xEnd[6], xEnd[5], xEnd[4], xEnd[3], xEnd[2], xEnd[1], xEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_91_ ), 
        .DX( {nn4467, nn4466, nn4465, nn4464, nn4463, nn4462, nn4461, nn4460, 
              nn4459, nn4458, nn4457, nn4456} ), 
        .SUM( {\inputctrl1_u41_XORCI_11|SUM_net , dummy_92_, dummy_93_, dummy_94_, 
              dummy_95_, dummy_96_, dummy_97_, dummy_98_, dummy_99_, dummy_100_, 
              dummy_101_, dummy_102_} )
      );
    CS_LUT4_PRIM ii4482 ( .DX(nn4482), .F0(yBgn[0]), .F1(\inputctrl1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_3223_), .F3(dummy_abc_3224_) );
      defparam ii4482.CONFIG_DATA = 16'h9999;
      defparam ii4482.PLACE_LOCATION = "NONE";
      defparam ii4482.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4483 ( .DX(nn4483), .F0(yBgn[1]), .F1(\inputctrl1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_3225_), .F3(dummy_abc_3226_) );
      defparam ii4483.CONFIG_DATA = 16'h9999;
      defparam ii4483.PLACE_LOCATION = "NONE";
      defparam ii4483.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4484 ( .DX(nn4484), .F0(yBgn[2]), .F1(\inputctrl1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_3227_), .F3(dummy_abc_3228_) );
      defparam ii4484.CONFIG_DATA = 16'h9999;
      defparam ii4484.PLACE_LOCATION = "NONE";
      defparam ii4484.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4485 ( .DX(nn4485), .F0(yBgn[3]), .F1(\inputctrl1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_3229_), .F3(dummy_abc_3230_) );
      defparam ii4485.CONFIG_DATA = 16'h9999;
      defparam ii4485.PLACE_LOCATION = "NONE";
      defparam ii4485.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4486 ( .DX(nn4486), .F0(yBgn[4]), .F1(\inputctrl1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_3231_), .F3(dummy_abc_3232_) );
      defparam ii4486.CONFIG_DATA = 16'h9999;
      defparam ii4486.PLACE_LOCATION = "NONE";
      defparam ii4486.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4487 ( .DX(nn4487), .F0(yBgn[5]), .F1(\inputctrl1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_3233_), .F3(dummy_abc_3234_) );
      defparam ii4487.CONFIG_DATA = 16'h9999;
      defparam ii4487.PLACE_LOCATION = "NONE";
      defparam ii4487.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4488 ( .DX(nn4488), .F0(yBgn[6]), .F1(\inputctrl1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_3235_), .F3(dummy_abc_3236_) );
      defparam ii4488.CONFIG_DATA = 16'h9999;
      defparam ii4488.PLACE_LOCATION = "NONE";
      defparam ii4488.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4489 ( .DX(nn4489), .F0(yBgn[7]), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_3237_), .F3(dummy_abc_3238_) );
      defparam ii4489.CONFIG_DATA = 16'h9999;
      defparam ii4489.PLACE_LOCATION = "NONE";
      defparam ii4489.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4490 ( .DX(nn4490), .F0(yBgn[8]), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_3239_), .F3(dummy_abc_3240_) );
      defparam ii4490.CONFIG_DATA = 16'h9999;
      defparam ii4490.PLACE_LOCATION = "NONE";
      defparam ii4490.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4491 ( .DX(nn4491), .F0(yBgn[9]), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_3241_), .F3(dummy_abc_3242_) );
      defparam ii4491.CONFIG_DATA = 16'h9999;
      defparam ii4491.PLACE_LOCATION = "NONE";
      defparam ii4491.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4492 ( .DX(nn4492), .F0(yBgn[10]), .F1(\inputctrl1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_3243_), .F3(dummy_abc_3244_) );
      defparam ii4492.CONFIG_DATA = 16'h9999;
      defparam ii4492.PLACE_LOCATION = "NONE";
      defparam ii4492.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4493 ( .DX(nn4493), .F0(dummy_abc_3245_), .F1(dummy_abc_3246_), .F2(dummy_abc_3247_), .F3(dummy_abc_3248_) );
      defparam ii4493.CONFIG_DATA = 16'hFFFF;
      defparam ii4493.PLACE_LOCATION = "NONE";
      defparam ii4493.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_83_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \inputctrl1_yAddress__reg[10]|Q_net , 
              \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net , 
              \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net , 
              \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net , 
              \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net , 
              \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_78_ ), 
        .DX( {nn4493, nn4492, nn4491, nn4490, nn4489, nn4488, nn4487, nn4486, 
              nn4485, nn4484, nn4483, nn4482} ), 
        .SUM( {\inputctrl1_u39_XORCI_11|SUM_net , dummy_79_, dummy_80_, dummy_81_, 
              dummy_82_, dummy_83_, dummy_84_, dummy_85_, dummy_86_, dummy_87_, 
              dummy_88_, dummy_89_} )
      );
    CS_LUT4_PRIM ii4508 ( .DX(nn4508), .F0(xBgn[0]), .F1(\inputctrl1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_3249_), .F3(dummy_abc_3250_) );
      defparam ii4508.CONFIG_DATA = 16'h9999;
      defparam ii4508.PLACE_LOCATION = "NONE";
      defparam ii4508.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4509 ( .DX(nn4509), .F0(xBgn[1]), .F1(\inputctrl1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_3251_), .F3(dummy_abc_3252_) );
      defparam ii4509.CONFIG_DATA = 16'h9999;
      defparam ii4509.PLACE_LOCATION = "NONE";
      defparam ii4509.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4510 ( .DX(nn4510), .F0(xBgn[2]), .F1(\inputctrl1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_3253_), .F3(dummy_abc_3254_) );
      defparam ii4510.CONFIG_DATA = 16'h9999;
      defparam ii4510.PLACE_LOCATION = "NONE";
      defparam ii4510.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4511 ( .DX(nn4511), .F0(xBgn[3]), .F1(\inputctrl1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_3255_), .F3(dummy_abc_3256_) );
      defparam ii4511.CONFIG_DATA = 16'h9999;
      defparam ii4511.PLACE_LOCATION = "NONE";
      defparam ii4511.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4512 ( .DX(nn4512), .F0(xBgn[4]), .F1(\inputctrl1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_3257_), .F3(dummy_abc_3258_) );
      defparam ii4512.CONFIG_DATA = 16'h9999;
      defparam ii4512.PLACE_LOCATION = "NONE";
      defparam ii4512.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4513 ( .DX(nn4513), .F0(xBgn[5]), .F1(\inputctrl1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_3259_), .F3(dummy_abc_3260_) );
      defparam ii4513.CONFIG_DATA = 16'h9999;
      defparam ii4513.PLACE_LOCATION = "NONE";
      defparam ii4513.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4514 ( .DX(nn4514), .F0(xBgn[6]), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_3261_), .F3(dummy_abc_3262_) );
      defparam ii4514.CONFIG_DATA = 16'h9999;
      defparam ii4514.PLACE_LOCATION = "NONE";
      defparam ii4514.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4515 ( .DX(nn4515), .F0(xBgn[7]), .F1(\inputctrl1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_3263_), .F3(dummy_abc_3264_) );
      defparam ii4515.CONFIG_DATA = 16'h9999;
      defparam ii4515.PLACE_LOCATION = "NONE";
      defparam ii4515.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4516 ( .DX(nn4516), .F0(xBgn[8]), .F1(\inputctrl1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_3265_), .F3(dummy_abc_3266_) );
      defparam ii4516.CONFIG_DATA = 16'h9999;
      defparam ii4516.PLACE_LOCATION = "NONE";
      defparam ii4516.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4517 ( .DX(nn4517), .F0(xBgn[9]), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_3267_), .F3(dummy_abc_3268_) );
      defparam ii4517.CONFIG_DATA = 16'h9999;
      defparam ii4517.PLACE_LOCATION = "NONE";
      defparam ii4517.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4518 ( .DX(nn4518), .F0(xBgn[10]), .F1(\inputctrl1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_3269_), .F3(dummy_abc_3270_) );
      defparam ii4518.CONFIG_DATA = 16'h9999;
      defparam ii4518.PLACE_LOCATION = "NONE";
      defparam ii4518.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4519 ( .DX(nn4519), .F0(dummy_abc_3271_), .F1(dummy_abc_3272_), .F2(dummy_abc_3273_), .F3(dummy_abc_3274_) );
      defparam ii4519.CONFIG_DATA = 16'hFFFF;
      defparam ii4519.PLACE_LOCATION = "NONE";
      defparam ii4519.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_82_ ( 
        .CA( {a_acc_en_cal1_u134_mac, \inputctrl1_xAddress__reg[10]|Q_net , 
              \inputctrl1_xAddress__reg[9]|Q_net , \inputctrl1_xAddress__reg[8]|Q_net , 
              \inputctrl1_xAddress__reg[7]|Q_net , \inputctrl1_xAddress__reg[6]|Q_net , 
              \inputctrl1_xAddress__reg[5]|Q_net , \inputctrl1_xAddress__reg[4]|Q_net , 
              \inputctrl1_xAddress__reg[3]|Q_net , \inputctrl1_xAddress__reg[2]|Q_net , 
              \inputctrl1_xAddress__reg[1]|Q_net , \inputctrl1_xAddress__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u134_mac ), 
        .CO( dummy_65_ ), 
        .DX( {nn4519, nn4518, nn4517, nn4516, nn4515, nn4514, nn4513, nn4512, 
              nn4511, nn4510, nn4509, nn4508} ), 
        .SUM( {\inputctrl1_u37_XORCI_11|SUM_net , dummy_66_, dummy_67_, dummy_68_, 
              dummy_69_, dummy_70_, dummy_71_, dummy_72_, dummy_73_, dummy_74_, 
              dummy_75_, dummy_76_} )
      );
    CS_LUT4_PRIM ii4534 ( .DX(nn4534), .F0(dInEn), .F1(dummy_91_), .F2(dummy_78_), .F3(dummy_65_) );
      defparam ii4534.CONFIG_DATA = 16'h8000;
      defparam ii4534.PLACE_LOCATION = "NONE";
      defparam ii4534.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4535 ( .DX(nn4535), .F0(\inputctrl1_xPreEn__reg|Q_net ), .F1(dummy_104_), .F2(nn4455), .F3(nn4534) );
      defparam ii4535.CONFIG_DATA = 16'hC800;
      defparam ii4535.PLACE_LOCATION = "NONE";
      defparam ii4535.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4536 ( .DX(nn4536), .F0(iHsyn), .F1(iVsyn), .F2(nn4422), .F3(nn4535) );
      defparam ii4536.CONFIG_DATA = 16'hEFEE;
      defparam ii4536.PLACE_LOCATION = "NONE";
      defparam ii4536.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4537 ( .DX(nn4537), .F0(dIn[10]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3275_) );
      defparam ii4537.CONFIG_DATA = 16'h0202;
      defparam ii4537.PLACE_LOCATION = "NONE";
      defparam ii4537.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4538 ( .DX(nn4538), .F0(dIn[11]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3276_) );
      defparam ii4538.CONFIG_DATA = 16'h0202;
      defparam ii4538.PLACE_LOCATION = "NONE";
      defparam ii4538.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4539 ( .DX(nn4539), .F0(dIn[12]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3277_) );
      defparam ii4539.CONFIG_DATA = 16'h0202;
      defparam ii4539.PLACE_LOCATION = "NONE";
      defparam ii4539.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4540 ( .DX(nn4540), .F0(dIn[13]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3278_) );
      defparam ii4540.CONFIG_DATA = 16'h0202;
      defparam ii4540.PLACE_LOCATION = "NONE";
      defparam ii4540.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4541 ( .DX(nn4541), .F0(dIn[14]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3279_) );
      defparam ii4541.CONFIG_DATA = 16'h0202;
      defparam ii4541.PLACE_LOCATION = "NONE";
      defparam ii4541.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4542 ( .DX(nn4542), .F0(dIn[15]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3280_) );
      defparam ii4542.CONFIG_DATA = 16'h0202;
      defparam ii4542.PLACE_LOCATION = "NONE";
      defparam ii4542.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4543 ( .DX(nn4543), .F0(dIn[1]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3281_) );
      defparam ii4543.CONFIG_DATA = 16'h0202;
      defparam ii4543.PLACE_LOCATION = "NONE";
      defparam ii4543.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4544 ( .DX(nn4544), .F0(dIn[2]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3282_) );
      defparam ii4544.CONFIG_DATA = 16'h0202;
      defparam ii4544.PLACE_LOCATION = "NONE";
      defparam ii4544.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4545 ( .DX(nn4545), .F0(dIn[3]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3283_) );
      defparam ii4545.CONFIG_DATA = 16'h0202;
      defparam ii4545.PLACE_LOCATION = "NONE";
      defparam ii4545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4546 ( .DX(nn4546), .F0(dIn[4]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3284_) );
      defparam ii4546.CONFIG_DATA = 16'h0202;
      defparam ii4546.PLACE_LOCATION = "NONE";
      defparam ii4546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4547 ( .DX(nn4547), .F0(dIn[5]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3285_) );
      defparam ii4547.CONFIG_DATA = 16'h0202;
      defparam ii4547.PLACE_LOCATION = "NONE";
      defparam ii4547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4548 ( .DX(nn4548), .F0(dIn[6]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3286_) );
      defparam ii4548.CONFIG_DATA = 16'h0202;
      defparam ii4548.PLACE_LOCATION = "NONE";
      defparam ii4548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4549 ( .DX(nn4549), .F0(dIn[7]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3287_) );
      defparam ii4549.CONFIG_DATA = 16'h0202;
      defparam ii4549.PLACE_LOCATION = "NONE";
      defparam ii4549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4550 ( .DX(nn4550), .F0(dIn[8]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3288_) );
      defparam ii4550.CONFIG_DATA = 16'h0202;
      defparam ii4550.PLACE_LOCATION = "NONE";
      defparam ii4550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4551 ( .DX(nn4551), .F0(dIn[9]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3289_) );
      defparam ii4551.CONFIG_DATA = 16'h0202;
      defparam ii4551.PLACE_LOCATION = "NONE";
      defparam ii4551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4552 ( .DX(nn4552), .F0(iHsyn), .F1(nn4422), .F2(dummy_abc_3290_), .F3(dummy_abc_3291_) );
      defparam ii4552.CONFIG_DATA = 16'h2222;
      defparam ii4552.PLACE_LOCATION = "NONE";
      defparam ii4552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4553 ( .DX(nn4553), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F3(dummy_abc_3292_) );
      defparam ii4553.CONFIG_DATA = 16'hEFEF;
      defparam ii4553.PLACE_LOCATION = "NONE";
      defparam ii4553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4554 ( .DX(nn4554), .F0(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F1(dummy_abc_3293_), .F2(dummy_abc_3294_), .F3(dummy_abc_3295_) );
      defparam ii4554.CONFIG_DATA = 16'h5555;
      defparam ii4554.PLACE_LOCATION = "NONE";
      defparam ii4554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4555 ( .DX(nn4555), .F0(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F1(dummy_abc_3296_), .F2(dummy_abc_3297_), .F3(dummy_abc_3298_) );
      defparam ii4555.CONFIG_DATA = 16'hAAAA;
      defparam ii4555.PLACE_LOCATION = "NONE";
      defparam ii4555.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4556 ( .DX(nn4556), .F0(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F1(dummy_abc_3299_), .F2(dummy_abc_3300_), .F3(dummy_abc_3301_) );
      defparam ii4556.CONFIG_DATA = 16'hAAAA;
      defparam ii4556.PLACE_LOCATION = "NONE";
      defparam ii4556.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4557 ( .DX(nn4557), .F0(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F1(dummy_abc_3302_), .F2(dummy_abc_3303_), .F3(dummy_abc_3304_) );
      defparam ii4557.CONFIG_DATA = 16'hAAAA;
      defparam ii4557.PLACE_LOCATION = "NONE";
      defparam ii4557.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4558 ( .DX(nn4558), .F0(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F1(dummy_abc_3305_), .F2(dummy_abc_3306_), .F3(dummy_abc_3307_) );
      defparam ii4558.CONFIG_DATA = 16'hAAAA;
      defparam ii4558.PLACE_LOCATION = "NONE";
      defparam ii4558.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4559 ( .DX(nn4559), .F0(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F1(dummy_abc_3308_), .F2(dummy_abc_3309_), .F3(dummy_abc_3310_) );
      defparam ii4559.CONFIG_DATA = 16'hAAAA;
      defparam ii4559.PLACE_LOCATION = "NONE";
      defparam ii4559.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4560 ( .DX(nn4560), .F0(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F1(dummy_abc_3311_), .F2(dummy_abc_3312_), .F3(dummy_abc_3313_) );
      defparam ii4560.CONFIG_DATA = 16'hAAAA;
      defparam ii4560.PLACE_LOCATION = "NONE";
      defparam ii4560.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4561 ( .DX(nn4561), .F0(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F1(dummy_abc_3314_), .F2(dummy_abc_3315_), .F3(dummy_abc_3316_) );
      defparam ii4561.CONFIG_DATA = 16'hAAAA;
      defparam ii4561.PLACE_LOCATION = "NONE";
      defparam ii4561.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4562 ( .DX(nn4562), .F0(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F1(dummy_abc_3317_), .F2(dummy_abc_3318_), .F3(dummy_abc_3319_) );
      defparam ii4562.CONFIG_DATA = 16'hAAAA;
      defparam ii4562.PLACE_LOCATION = "NONE";
      defparam ii4562.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4563 ( .DX(nn4563), .F0(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F1(dummy_abc_3320_), .F2(dummy_abc_3321_), .F3(dummy_abc_3322_) );
      defparam ii4563.CONFIG_DATA = 16'hAAAA;
      defparam ii4563.PLACE_LOCATION = "NONE";
      defparam ii4563.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4564 ( .DX(nn4564), .F0(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F1(dummy_abc_3323_), .F2(dummy_abc_3324_), .F3(dummy_abc_3325_) );
      defparam ii4564.CONFIG_DATA = 16'hAAAA;
      defparam ii4564.PLACE_LOCATION = "NONE";
      defparam ii4564.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_81_ ( 
        .CA( {\inputctrl1_ramWrtAddr__reg[10]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[9]|Q_net , \inputctrl1_ramWrtAddr__reg[8]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[7]|Q_net , \inputctrl1_ramWrtAddr__reg[6]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[5]|Q_net , \inputctrl1_ramWrtAddr__reg[4]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[3]|Q_net , \inputctrl1_ramWrtAddr__reg[2]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[1]|Q_net , \inputctrl1_ramWrtAddr__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_20_ ), 
        .DX( {nn4564, nn4563, nn4562, nn4561, nn4560, nn4559, nn4558, nn4557, 
              nn4556, nn4555, nn4554} ), 
        .SUM( {\inputctrl1_u112_XORCI_10|SUM_net , 
              \inputctrl1_u112_XORCI_9|SUM_net , \inputctrl1_u112_XORCI_8|SUM_net , 
              \inputctrl1_u112_XORCI_7|SUM_net , \inputctrl1_u112_XORCI_6|SUM_net , 
              \inputctrl1_u112_XORCI_5|SUM_net , \inputctrl1_u112_XORCI_4|SUM_net , 
              \inputctrl1_u112_XORCI_3|SUM_net , \inputctrl1_u112_XORCI_2|SUM_net , 
              \inputctrl1_u112_XORCI_1|SUM_net , \inputctrl1_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4578 ( .DX(nn4578), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_10|SUM_net ), .F3(dummy_abc_3326_) );
      defparam ii4578.CONFIG_DATA = 16'hFEFE;
      defparam ii4578.PLACE_LOCATION = "NONE";
      defparam ii4578.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4579 ( .DX(nn4579), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_1|SUM_net ), .F3(dummy_abc_3327_) );
      defparam ii4579.CONFIG_DATA = 16'hFEFE;
      defparam ii4579.PLACE_LOCATION = "NONE";
      defparam ii4579.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4580 ( .DX(nn4580), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_2|SUM_net ), .F3(dummy_abc_3328_) );
      defparam ii4580.CONFIG_DATA = 16'hFEFE;
      defparam ii4580.PLACE_LOCATION = "NONE";
      defparam ii4580.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4581 ( .DX(nn4581), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_3|SUM_net ), .F3(dummy_abc_3329_) );
      defparam ii4581.CONFIG_DATA = 16'hFEFE;
      defparam ii4581.PLACE_LOCATION = "NONE";
      defparam ii4581.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4582 ( .DX(nn4582), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_4|SUM_net ), .F3(dummy_abc_3330_) );
      defparam ii4582.CONFIG_DATA = 16'hFEFE;
      defparam ii4582.PLACE_LOCATION = "NONE";
      defparam ii4582.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4583 ( .DX(nn4583), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_5|SUM_net ), .F3(dummy_abc_3331_) );
      defparam ii4583.CONFIG_DATA = 16'hFEFE;
      defparam ii4583.PLACE_LOCATION = "NONE";
      defparam ii4583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4584 ( .DX(nn4584), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_6|SUM_net ), .F3(dummy_abc_3332_) );
      defparam ii4584.CONFIG_DATA = 16'hFEFE;
      defparam ii4584.PLACE_LOCATION = "NONE";
      defparam ii4584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4585 ( .DX(nn4585), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_7|SUM_net ), .F3(dummy_abc_3333_) );
      defparam ii4585.CONFIG_DATA = 16'hFEFE;
      defparam ii4585.PLACE_LOCATION = "NONE";
      defparam ii4585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4586 ( .DX(nn4586), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_8|SUM_net ), .F3(dummy_abc_3334_) );
      defparam ii4586.CONFIG_DATA = 16'hFEFE;
      defparam ii4586.PLACE_LOCATION = "NONE";
      defparam ii4586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4587 ( .DX(nn4587), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_9|SUM_net ), .F3(dummy_abc_3335_) );
      defparam ii4587.CONFIG_DATA = 16'hFEFE;
      defparam ii4587.PLACE_LOCATION = "NONE";
      defparam ii4587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4588 ( .DX(nn4588), .F0(iHsyn), .F1(iVsyn), .F2(nn4422), .F3(nn4535) );
      defparam ii4588.CONFIG_DATA = 16'h0100;
      defparam ii4588.PLACE_LOCATION = "NONE";
      defparam ii4588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4589 ( .DX(nn4589), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_3336_), .F2(dummy_abc_3337_), .F3(dummy_abc_3338_) );
      defparam ii4589.CONFIG_DATA = 16'h5555;
      defparam ii4589.PLACE_LOCATION = "NONE";
      defparam ii4589.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4590 ( .DX(nn4590), .F0(iHsyn), .F1(iVsyn), .F2(rst), .F3(\coefcal1_inEn__reg|Q_net ) );
      defparam ii4590.CONFIG_DATA = 16'hFEF0;
      defparam ii4590.PLACE_LOCATION = "NONE";
      defparam ii4590.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4591 ( .DX(nn4591), .F0(dInEn), .F1(\coefcal1_inEn__reg|Q_net ), .F2(dummy_abc_3339_), .F3(dummy_abc_3340_) );
      defparam ii4591.CONFIG_DATA = 16'h8888;
      defparam ii4591.PLACE_LOCATION = "NONE";
      defparam ii4591.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4592 ( .DX(nn4592), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_3341_), .F2(dummy_abc_3342_), .F3(dummy_abc_3343_) );
      defparam ii4592.CONFIG_DATA = 16'h5555;
      defparam ii4592.PLACE_LOCATION = "NONE";
      defparam ii4592.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4593 ( .DX(nn4593), .F0(\inputctrl1_xAddress__reg[1]|Q_net ), .F1(dummy_abc_3344_), .F2(dummy_abc_3345_), .F3(dummy_abc_3346_) );
      defparam ii4593.CONFIG_DATA = 16'hAAAA;
      defparam ii4593.PLACE_LOCATION = "NONE";
      defparam ii4593.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4594 ( .DX(nn4594), .F0(\inputctrl1_xAddress__reg[2]|Q_net ), .F1(dummy_abc_3347_), .F2(dummy_abc_3348_), .F3(dummy_abc_3349_) );
      defparam ii4594.CONFIG_DATA = 16'hAAAA;
      defparam ii4594.PLACE_LOCATION = "NONE";
      defparam ii4594.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4595 ( .DX(nn4595), .F0(\inputctrl1_xAddress__reg[3]|Q_net ), .F1(dummy_abc_3350_), .F2(dummy_abc_3351_), .F3(dummy_abc_3352_) );
      defparam ii4595.CONFIG_DATA = 16'hAAAA;
      defparam ii4595.PLACE_LOCATION = "NONE";
      defparam ii4595.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4596 ( .DX(nn4596), .F0(\inputctrl1_xAddress__reg[4]|Q_net ), .F1(dummy_abc_3353_), .F2(dummy_abc_3354_), .F3(dummy_abc_3355_) );
      defparam ii4596.CONFIG_DATA = 16'hAAAA;
      defparam ii4596.PLACE_LOCATION = "NONE";
      defparam ii4596.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4597 ( .DX(nn4597), .F0(\inputctrl1_xAddress__reg[5]|Q_net ), .F1(dummy_abc_3356_), .F2(dummy_abc_3357_), .F3(dummy_abc_3358_) );
      defparam ii4597.CONFIG_DATA = 16'hAAAA;
      defparam ii4597.PLACE_LOCATION = "NONE";
      defparam ii4597.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4598 ( .DX(nn4598), .F0(\inputctrl1_xAddress__reg[6]|Q_net ), .F1(dummy_abc_3359_), .F2(dummy_abc_3360_), .F3(dummy_abc_3361_) );
      defparam ii4598.CONFIG_DATA = 16'hAAAA;
      defparam ii4598.PLACE_LOCATION = "NONE";
      defparam ii4598.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4599 ( .DX(nn4599), .F0(\inputctrl1_xAddress__reg[7]|Q_net ), .F1(dummy_abc_3362_), .F2(dummy_abc_3363_), .F3(dummy_abc_3364_) );
      defparam ii4599.CONFIG_DATA = 16'hAAAA;
      defparam ii4599.PLACE_LOCATION = "NONE";
      defparam ii4599.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4600 ( .DX(nn4600), .F0(\inputctrl1_xAddress__reg[8]|Q_net ), .F1(dummy_abc_3365_), .F2(dummy_abc_3366_), .F3(dummy_abc_3367_) );
      defparam ii4600.CONFIG_DATA = 16'hAAAA;
      defparam ii4600.PLACE_LOCATION = "NONE";
      defparam ii4600.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4601 ( .DX(nn4601), .F0(\inputctrl1_xAddress__reg[9]|Q_net ), .F1(dummy_abc_3368_), .F2(dummy_abc_3369_), .F3(dummy_abc_3370_) );
      defparam ii4601.CONFIG_DATA = 16'hAAAA;
      defparam ii4601.PLACE_LOCATION = "NONE";
      defparam ii4601.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4602 ( .DX(nn4602), .F0(\inputctrl1_xAddress__reg[10]|Q_net ), .F1(dummy_abc_3371_), .F2(dummy_abc_3372_), .F3(dummy_abc_3373_) );
      defparam ii4602.CONFIG_DATA = 16'hAAAA;
      defparam ii4602.PLACE_LOCATION = "NONE";
      defparam ii4602.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_79_ ( 
        .CA( {\inputctrl1_xAddress__reg[10]|Q_net , 
              \inputctrl1_xAddress__reg[9]|Q_net , \inputctrl1_xAddress__reg[8]|Q_net , 
              \inputctrl1_xAddress__reg[7]|Q_net , \inputctrl1_xAddress__reg[6]|Q_net , 
              \inputctrl1_xAddress__reg[5]|Q_net , \inputctrl1_xAddress__reg[4]|Q_net , 
              \inputctrl1_xAddress__reg[3]|Q_net , \inputctrl1_xAddress__reg[2]|Q_net , 
              \inputctrl1_xAddress__reg[1]|Q_net , \inputctrl1_xAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_18_ ), 
        .DX( {nn4602, nn4601, nn4600, nn4599, nn4598, nn4597, nn4596, nn4595, 
              nn4594, nn4593, nn4592} ), 
        .SUM( {\inputctrl1_u110_XORCI_10|SUM_net , 
              \inputctrl1_u110_XORCI_9|SUM_net , \inputctrl1_u110_XORCI_8|SUM_net , 
              \inputctrl1_u110_XORCI_7|SUM_net , \inputctrl1_u110_XORCI_6|SUM_net , 
              \inputctrl1_u110_XORCI_5|SUM_net , \inputctrl1_u110_XORCI_4|SUM_net , 
              \inputctrl1_u110_XORCI_3|SUM_net , \inputctrl1_u110_XORCI_2|SUM_net , 
              \inputctrl1_u110_XORCI_1|SUM_net , \inputctrl1_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4616 ( .DX(nn4616), .F0(\coefcal1_u61_XORCI_6|SUM_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_65_), .F3(dummy_abc_3374_) );
      defparam ii4616.CONFIG_DATA = 16'hE0E0;
      defparam ii4616.PLACE_LOCATION = "NONE";
      defparam ii4616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4617 ( .DX(nn4617), .F0(\inputctrl1_xCal__reg[0]|Q_net ), .F1(nn4025), .F2(nn4616), .F3(dummy_abc_3375_) );
      defparam ii4617.CONFIG_DATA = 16'h6A6A;
      defparam ii4617.PLACE_LOCATION = "NONE";
      defparam ii4617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4618 ( .DX(nn4618), .F0(nn4455), .F1(nn4591), .F2(dummy_abc_3376_), .F3(dummy_abc_3377_) );
      defparam ii4618.CONFIG_DATA = 16'h8888;
      defparam ii4618.PLACE_LOCATION = "NONE";
      defparam ii4618.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4619 ( .DX(nn4619), .F0(\inputctrl1_xCal__reg[0]|Q_net ), .F1(nn4025), .F2(nn4616), .F3(dummy_abc_3378_) );
      defparam ii4619.CONFIG_DATA = 16'h6A6A;
      defparam ii4619.PLACE_LOCATION = "NONE";
      defparam ii4619.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4620 ( .DX(nn4620), .F0(\inputctrl1_xCal__reg[1]|Q_net ), .F1(\coefcal1_u61_XORCI_1|SUM_net ), .F2(nn4616), .F3(dummy_abc_3379_) );
      defparam ii4620.CONFIG_DATA = 16'h6A6A;
      defparam ii4620.PLACE_LOCATION = "NONE";
      defparam ii4620.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4621 ( .DX(nn4621), .F0(\inputctrl1_xCal__reg[2]|Q_net ), .F1(\coefcal1_u61_XORCI_2|SUM_net ), .F2(nn4616), .F3(dummy_abc_3380_) );
      defparam ii4621.CONFIG_DATA = 16'h6A6A;
      defparam ii4621.PLACE_LOCATION = "NONE";
      defparam ii4621.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4622 ( .DX(nn4622), .F0(\inputctrl1_xCal__reg[3]|Q_net ), .F1(\coefcal1_u61_XORCI_3|SUM_net ), .F2(nn4616), .F3(dummy_abc_3381_) );
      defparam ii4622.CONFIG_DATA = 16'h6A6A;
      defparam ii4622.PLACE_LOCATION = "NONE";
      defparam ii4622.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4623 ( .DX(nn4623), .F0(\inputctrl1_xCal__reg[4]|Q_net ), .F1(\coefcal1_u61_XORCI_4|SUM_net ), .F2(nn4616), .F3(dummy_abc_3382_) );
      defparam ii4623.CONFIG_DATA = 16'h6A6A;
      defparam ii4623.PLACE_LOCATION = "NONE";
      defparam ii4623.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4624 ( .DX(nn4624), .F0(\inputctrl1_xCal__reg[5]|Q_net ), .F1(\coefcal1_u61_XORCI_5|SUM_net ), .F2(nn4616), .F3(dummy_abc_3383_) );
      defparam ii4624.CONFIG_DATA = 16'h6A6A;
      defparam ii4624.PLACE_LOCATION = "NONE";
      defparam ii4624.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4625 ( .DX(nn4625), .F0(\inputctrl1_xCal__reg[6]|Q_net ), .F1(\coefcal1_u61_XORCI_6|SUM_net ), .F2(nn4616), .F3(dummy_abc_3384_) );
      defparam ii4625.CONFIG_DATA = 16'h6565;
      defparam ii4625.PLACE_LOCATION = "NONE";
      defparam ii4625.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4626 ( .DX(nn4626), .F0(\inputctrl1_xCal__reg[7]|Q_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_65_), .F3(dummy_abc_3385_) );
      defparam ii4626.CONFIG_DATA = 16'h6A6A;
      defparam ii4626.PLACE_LOCATION = "NONE";
      defparam ii4626.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4627 ( .DX(nn4627), .F0(\inputctrl1_xCal__reg[8]|Q_net ), .F1(dummy_abc_3386_), .F2(dummy_abc_3387_), .F3(dummy_abc_3388_) );
      defparam ii4627.CONFIG_DATA = 16'hAAAA;
      defparam ii4627.PLACE_LOCATION = "NONE";
      defparam ii4627.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4628 ( .DX(nn4628), .F0(\inputctrl1_xCal__reg[9]|Q_net ), .F1(dummy_abc_3389_), .F2(dummy_abc_3390_), .F3(dummy_abc_3391_) );
      defparam ii4628.CONFIG_DATA = 16'hAAAA;
      defparam ii4628.PLACE_LOCATION = "NONE";
      defparam ii4628.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4629 ( .DX(nn4629), .F0(\inputctrl1_xCal__reg[10]|Q_net ), .F1(dummy_abc_3392_), .F2(dummy_abc_3393_), .F3(dummy_abc_3394_) );
      defparam ii4629.CONFIG_DATA = 16'hAAAA;
      defparam ii4629.PLACE_LOCATION = "NONE";
      defparam ii4629.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4630 ( .DX(nn4630), .F0(\inputctrl1_xCal__reg[11]|Q_net ), .F1(dummy_abc_3395_), .F2(dummy_abc_3396_), .F3(dummy_abc_3397_) );
      defparam ii4630.CONFIG_DATA = 16'hAAAA;
      defparam ii4630.PLACE_LOCATION = "NONE";
      defparam ii4630.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4631 ( .DX(nn4631), .F0(\inputctrl1_xCal__reg[12]|Q_net ), .F1(dummy_abc_3398_), .F2(dummy_abc_3399_), .F3(dummy_abc_3400_) );
      defparam ii4631.CONFIG_DATA = 16'hAAAA;
      defparam ii4631.PLACE_LOCATION = "NONE";
      defparam ii4631.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4632 ( .DX(nn4632), .F0(\inputctrl1_xCal__reg[13]|Q_net ), .F1(dummy_abc_3401_), .F2(dummy_abc_3402_), .F3(dummy_abc_3403_) );
      defparam ii4632.CONFIG_DATA = 16'hAAAA;
      defparam ii4632.PLACE_LOCATION = "NONE";
      defparam ii4632.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4633 ( .DX(nn4633), .F0(\inputctrl1_xCal__reg[14]|Q_net ), .F1(dummy_abc_3404_), .F2(dummy_abc_3405_), .F3(dummy_abc_3406_) );
      defparam ii4633.CONFIG_DATA = 16'hAAAA;
      defparam ii4633.PLACE_LOCATION = "NONE";
      defparam ii4633.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4634 ( .DX(nn4634), .F0(\inputctrl1_xCal__reg[15]|Q_net ), .F1(dummy_abc_3407_), .F2(dummy_abc_3408_), .F3(dummy_abc_3409_) );
      defparam ii4634.CONFIG_DATA = 16'hAAAA;
      defparam ii4634.PLACE_LOCATION = "NONE";
      defparam ii4634.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4635 ( .DX(nn4635), .F0(\inputctrl1_xCal__reg[16]|Q_net ), .F1(dummy_abc_3410_), .F2(dummy_abc_3411_), .F3(dummy_abc_3412_) );
      defparam ii4635.CONFIG_DATA = 16'hAAAA;
      defparam ii4635.PLACE_LOCATION = "NONE";
      defparam ii4635.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_77_ ( 
        .CA( {\inputctrl1_xCal__reg[16]|Q_net , \inputctrl1_xCal__reg[15]|Q_net , 
              \inputctrl1_xCal__reg[14]|Q_net , \inputctrl1_xCal__reg[13]|Q_net , 
              \inputctrl1_xCal__reg[12]|Q_net , \inputctrl1_xCal__reg[11]|Q_net , 
              \inputctrl1_xCal__reg[10]|Q_net , \inputctrl1_xCal__reg[9]|Q_net , 
              \inputctrl1_xCal__reg[8]|Q_net , \inputctrl1_xCal__reg[7]|Q_net , 
              \inputctrl1_xCal__reg[6]|Q_net , \inputctrl1_xCal__reg[5]|Q_net , 
              \inputctrl1_xCal__reg[4]|Q_net , \inputctrl1_xCal__reg[3]|Q_net , 
              \inputctrl1_xCal__reg[2]|Q_net , \inputctrl1_xCal__reg[1]|Q_net , 
              \inputctrl1_xCal__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_198_ ), 
        .DX( {nn4635, nn4634, nn4633, nn4632, nn4631, nn4630, nn4629, nn4628, 
              nn4627, nn4626, nn4625, nn4624, nn4623, nn4622, nn4621, nn4620, 
              nn4619} ), 
        .SUM( {\inputctrl1_u108_XORCI_16|SUM_net , 
              \inputctrl1_u108_XORCI_15|SUM_net , \inputctrl1_u108_XORCI_14|SUM_net , 
              \inputctrl1_u108_XORCI_13|SUM_net , \inputctrl1_u108_XORCI_12|SUM_net , 
              \inputctrl1_u108_XORCI_11|SUM_net , \inputctrl1_u108_XORCI_10|SUM_net , 
              \inputctrl1_u108_XORCI_9|SUM_net , \inputctrl1_u108_XORCI_8|SUM_net , 
              \inputctrl1_u108_XORCI_7|SUM_net , \inputctrl1_u108_XORCI_6|SUM_net , 
              \inputctrl1_u108_XORCI_5|SUM_net , \inputctrl1_u108_XORCI_4|SUM_net , 
              \inputctrl1_u108_XORCI_3|SUM_net , \inputctrl1_u108_XORCI_2|SUM_net , 
              \inputctrl1_u108_XORCI_1|SUM_net , \inputctrl1_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4655 ( .DX(nn4655), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_3413_), .F2(dummy_abc_3414_), .F3(dummy_abc_3415_) );
      defparam ii4655.CONFIG_DATA = 16'h5555;
      defparam ii4655.PLACE_LOCATION = "NONE";
      defparam ii4655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4656 ( .DX(nn4656), .F0(iVsyn), .F1(rst), .F2(\coefcal1_inEn__reg|Q_net ), .F3(dummy_abc_3416_) );
      defparam ii4656.CONFIG_DATA = 16'hECEC;
      defparam ii4656.PLACE_LOCATION = "NONE";
      defparam ii4656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4657 ( .DX(nn4657), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_3417_), .F2(dummy_abc_3418_), .F3(dummy_abc_3419_) );
      defparam ii4657.CONFIG_DATA = 16'h5555;
      defparam ii4657.PLACE_LOCATION = "NONE";
      defparam ii4657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4658 ( .DX(nn4658), .F0(\inputctrl1_yAddress__reg[1]|Q_net ), .F1(dummy_abc_3420_), .F2(dummy_abc_3421_), .F3(dummy_abc_3422_) );
      defparam ii4658.CONFIG_DATA = 16'hAAAA;
      defparam ii4658.PLACE_LOCATION = "NONE";
      defparam ii4658.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4659 ( .DX(nn4659), .F0(\inputctrl1_yAddress__reg[2]|Q_net ), .F1(dummy_abc_3423_), .F2(dummy_abc_3424_), .F3(dummy_abc_3425_) );
      defparam ii4659.CONFIG_DATA = 16'hAAAA;
      defparam ii4659.PLACE_LOCATION = "NONE";
      defparam ii4659.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4660 ( .DX(nn4660), .F0(\inputctrl1_yAddress__reg[3]|Q_net ), .F1(dummy_abc_3426_), .F2(dummy_abc_3427_), .F3(dummy_abc_3428_) );
      defparam ii4660.CONFIG_DATA = 16'hAAAA;
      defparam ii4660.PLACE_LOCATION = "NONE";
      defparam ii4660.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4661 ( .DX(nn4661), .F0(\inputctrl1_yAddress__reg[4]|Q_net ), .F1(dummy_abc_3429_), .F2(dummy_abc_3430_), .F3(dummy_abc_3431_) );
      defparam ii4661.CONFIG_DATA = 16'hAAAA;
      defparam ii4661.PLACE_LOCATION = "NONE";
      defparam ii4661.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4662 ( .DX(nn4662), .F0(\inputctrl1_yAddress__reg[5]|Q_net ), .F1(dummy_abc_3432_), .F2(dummy_abc_3433_), .F3(dummy_abc_3434_) );
      defparam ii4662.CONFIG_DATA = 16'hAAAA;
      defparam ii4662.PLACE_LOCATION = "NONE";
      defparam ii4662.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4663 ( .DX(nn4663), .F0(\inputctrl1_yAddress__reg[6]|Q_net ), .F1(dummy_abc_3435_), .F2(dummy_abc_3436_), .F3(dummy_abc_3437_) );
      defparam ii4663.CONFIG_DATA = 16'hAAAA;
      defparam ii4663.PLACE_LOCATION = "NONE";
      defparam ii4663.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4664 ( .DX(nn4664), .F0(\inputctrl1_yAddress__reg[7]|Q_net ), .F1(dummy_abc_3438_), .F2(dummy_abc_3439_), .F3(dummy_abc_3440_) );
      defparam ii4664.CONFIG_DATA = 16'hAAAA;
      defparam ii4664.PLACE_LOCATION = "NONE";
      defparam ii4664.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4665 ( .DX(nn4665), .F0(\inputctrl1_yAddress__reg[8]|Q_net ), .F1(dummy_abc_3441_), .F2(dummy_abc_3442_), .F3(dummy_abc_3443_) );
      defparam ii4665.CONFIG_DATA = 16'hAAAA;
      defparam ii4665.PLACE_LOCATION = "NONE";
      defparam ii4665.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4666 ( .DX(nn4666), .F0(\inputctrl1_yAddress__reg[9]|Q_net ), .F1(dummy_abc_3444_), .F2(dummy_abc_3445_), .F3(dummy_abc_3446_) );
      defparam ii4666.CONFIG_DATA = 16'hAAAA;
      defparam ii4666.PLACE_LOCATION = "NONE";
      defparam ii4666.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4667 ( .DX(nn4667), .F0(\inputctrl1_yAddress__reg[10]|Q_net ), .F1(dummy_abc_3447_), .F2(dummy_abc_3448_), .F3(dummy_abc_3449_) );
      defparam ii4667.CONFIG_DATA = 16'hAAAA;
      defparam ii4667.PLACE_LOCATION = "NONE";
      defparam ii4667.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_80_ ( 
        .CA( {\inputctrl1_yAddress__reg[10]|Q_net , 
              \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net , 
              \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net , 
              \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net , 
              \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net , 
              \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_19_ ), 
        .DX( {nn4667, nn4666, nn4665, nn4664, nn4663, nn4662, nn4661, nn4660, 
              nn4659, nn4658, nn4657} ), 
        .SUM( {\inputctrl1_u111_XORCI_10|SUM_net , 
              \inputctrl1_u111_XORCI_9|SUM_net , \inputctrl1_u111_XORCI_8|SUM_net , 
              \inputctrl1_u111_XORCI_7|SUM_net , \inputctrl1_u111_XORCI_6|SUM_net , 
              \inputctrl1_u111_XORCI_5|SUM_net , \inputctrl1_u111_XORCI_4|SUM_net , 
              \inputctrl1_u111_XORCI_3|SUM_net , \inputctrl1_u111_XORCI_2|SUM_net , 
              \inputctrl1_u111_XORCI_1|SUM_net , \inputctrl1_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4681 ( .DX(nn4681), .F0(rst), .F1(dummy_526_), .F2(nn2644), .F3(dummy_abc_3450_) );
      defparam ii4681.CONFIG_DATA = 16'hFBFB;
      defparam ii4681.PLACE_LOCATION = "NONE";
      defparam ii4681.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4682 ( .DX(nn4682), .F0(\coefcal1_u62_XORCI_6|SUM_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_78_), .F3(dummy_abc_3451_) );
      defparam ii4682.CONFIG_DATA = 16'hE0E0;
      defparam ii4682.PLACE_LOCATION = "NONE";
      defparam ii4682.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4683 ( .DX(nn4683), .F0(\inputctrl1_yCal__reg[0]|Q_net ), .F1(nn4681), .F2(nn4682), .F3(dummy_abc_3452_) );
      defparam ii4683.CONFIG_DATA = 16'h6A6A;
      defparam ii4683.PLACE_LOCATION = "NONE";
      defparam ii4683.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4684 ( .DX(nn4684), .F0(iHsyn), .F1(nn4421), .F2(dummy_abc_3453_), .F3(dummy_abc_3454_) );
      defparam ii4684.CONFIG_DATA = 16'h8888;
      defparam ii4684.PLACE_LOCATION = "NONE";
      defparam ii4684.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4685 ( .DX(nn4685), .F0(\inputctrl1_yCal__reg[0]|Q_net ), .F1(nn4681), .F2(nn4682), .F3(dummy_abc_3455_) );
      defparam ii4685.CONFIG_DATA = 16'h6A6A;
      defparam ii4685.PLACE_LOCATION = "NONE";
      defparam ii4685.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4686 ( .DX(nn4686), .F0(\inputctrl1_yCal__reg[1]|Q_net ), .F1(\coefcal1_u62_XORCI_1|SUM_net ), .F2(nn4682), .F3(dummy_abc_3456_) );
      defparam ii4686.CONFIG_DATA = 16'h6A6A;
      defparam ii4686.PLACE_LOCATION = "NONE";
      defparam ii4686.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4687 ( .DX(nn4687), .F0(\inputctrl1_yCal__reg[2]|Q_net ), .F1(\coefcal1_u62_XORCI_2|SUM_net ), .F2(nn4682), .F3(dummy_abc_3457_) );
      defparam ii4687.CONFIG_DATA = 16'h6A6A;
      defparam ii4687.PLACE_LOCATION = "NONE";
      defparam ii4687.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4688 ( .DX(nn4688), .F0(\inputctrl1_yCal__reg[3]|Q_net ), .F1(\coefcal1_u62_XORCI_3|SUM_net ), .F2(nn4682), .F3(dummy_abc_3458_) );
      defparam ii4688.CONFIG_DATA = 16'h6A6A;
      defparam ii4688.PLACE_LOCATION = "NONE";
      defparam ii4688.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4689 ( .DX(nn4689), .F0(\inputctrl1_yCal__reg[4]|Q_net ), .F1(\coefcal1_u62_XORCI_4|SUM_net ), .F2(nn4682), .F3(dummy_abc_3459_) );
      defparam ii4689.CONFIG_DATA = 16'h6A6A;
      defparam ii4689.PLACE_LOCATION = "NONE";
      defparam ii4689.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4690 ( .DX(nn4690), .F0(\inputctrl1_yCal__reg[5]|Q_net ), .F1(\coefcal1_u62_XORCI_5|SUM_net ), .F2(nn4682), .F3(dummy_abc_3460_) );
      defparam ii4690.CONFIG_DATA = 16'h6A6A;
      defparam ii4690.PLACE_LOCATION = "NONE";
      defparam ii4690.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4691 ( .DX(nn4691), .F0(\inputctrl1_yCal__reg[6]|Q_net ), .F1(\coefcal1_u62_XORCI_6|SUM_net ), .F2(nn4682), .F3(dummy_abc_3461_) );
      defparam ii4691.CONFIG_DATA = 16'h6565;
      defparam ii4691.PLACE_LOCATION = "NONE";
      defparam ii4691.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4692 ( .DX(nn4692), .F0(\inputctrl1_yCal__reg[7]|Q_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_78_), .F3(dummy_abc_3462_) );
      defparam ii4692.CONFIG_DATA = 16'h6A6A;
      defparam ii4692.PLACE_LOCATION = "NONE";
      defparam ii4692.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4693 ( .DX(nn4693), .F0(\inputctrl1_yCal__reg[8]|Q_net ), .F1(dummy_abc_3463_), .F2(dummy_abc_3464_), .F3(dummy_abc_3465_) );
      defparam ii4693.CONFIG_DATA = 16'hAAAA;
      defparam ii4693.PLACE_LOCATION = "NONE";
      defparam ii4693.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4694 ( .DX(nn4694), .F0(\inputctrl1_yCal__reg[9]|Q_net ), .F1(dummy_abc_3466_), .F2(dummy_abc_3467_), .F3(dummy_abc_3468_) );
      defparam ii4694.CONFIG_DATA = 16'hAAAA;
      defparam ii4694.PLACE_LOCATION = "NONE";
      defparam ii4694.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4695 ( .DX(nn4695), .F0(\inputctrl1_yCal__reg[10]|Q_net ), .F1(dummy_abc_3469_), .F2(dummy_abc_3470_), .F3(dummy_abc_3471_) );
      defparam ii4695.CONFIG_DATA = 16'hAAAA;
      defparam ii4695.PLACE_LOCATION = "NONE";
      defparam ii4695.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4696 ( .DX(nn4696), .F0(\inputctrl1_yCal__reg[11]|Q_net ), .F1(dummy_abc_3472_), .F2(dummy_abc_3473_), .F3(dummy_abc_3474_) );
      defparam ii4696.CONFIG_DATA = 16'hAAAA;
      defparam ii4696.PLACE_LOCATION = "NONE";
      defparam ii4696.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4697 ( .DX(nn4697), .F0(\inputctrl1_yCal__reg[12]|Q_net ), .F1(dummy_abc_3475_), .F2(dummy_abc_3476_), .F3(dummy_abc_3477_) );
      defparam ii4697.CONFIG_DATA = 16'hAAAA;
      defparam ii4697.PLACE_LOCATION = "NONE";
      defparam ii4697.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4698 ( .DX(nn4698), .F0(\inputctrl1_yCal__reg[13]|Q_net ), .F1(dummy_abc_3478_), .F2(dummy_abc_3479_), .F3(dummy_abc_3480_) );
      defparam ii4698.CONFIG_DATA = 16'hAAAA;
      defparam ii4698.PLACE_LOCATION = "NONE";
      defparam ii4698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4699 ( .DX(nn4699), .F0(\inputctrl1_yCal__reg[14]|Q_net ), .F1(dummy_abc_3481_), .F2(dummy_abc_3482_), .F3(dummy_abc_3483_) );
      defparam ii4699.CONFIG_DATA = 16'hAAAA;
      defparam ii4699.PLACE_LOCATION = "NONE";
      defparam ii4699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4700 ( .DX(nn4700), .F0(\inputctrl1_yCal__reg[15]|Q_net ), .F1(dummy_abc_3484_), .F2(dummy_abc_3485_), .F3(dummy_abc_3486_) );
      defparam ii4700.CONFIG_DATA = 16'hAAAA;
      defparam ii4700.PLACE_LOCATION = "NONE";
      defparam ii4700.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4701 ( .DX(nn4701), .F0(\inputctrl1_yCal__reg[16]|Q_net ), .F1(dummy_abc_3487_), .F2(dummy_abc_3488_), .F3(dummy_abc_3489_) );
      defparam ii4701.CONFIG_DATA = 16'hAAAA;
      defparam ii4701.PLACE_LOCATION = "NONE";
      defparam ii4701.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_78_ ( 
        .CA( {\inputctrl1_yCal__reg[16]|Q_net , \inputctrl1_yCal__reg[15]|Q_net , 
              \inputctrl1_yCal__reg[14]|Q_net , \inputctrl1_yCal__reg[13]|Q_net , 
              \inputctrl1_yCal__reg[12]|Q_net , \inputctrl1_yCal__reg[11]|Q_net , 
              \inputctrl1_yCal__reg[10]|Q_net , \inputctrl1_yCal__reg[9]|Q_net , 
              \inputctrl1_yCal__reg[8]|Q_net , \inputctrl1_yCal__reg[7]|Q_net , 
              \inputctrl1_yCal__reg[6]|Q_net , \inputctrl1_yCal__reg[5]|Q_net , 
              \inputctrl1_yCal__reg[4]|Q_net , \inputctrl1_yCal__reg[3]|Q_net , 
              \inputctrl1_yCal__reg[2]|Q_net , \inputctrl1_yCal__reg[1]|Q_net , 
              \inputctrl1_yCal__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u134_mac ), 
        .CO( dummy_199_ ), 
        .DX( {nn4701, nn4700, nn4699, nn4698, nn4697, nn4696, nn4695, nn4694, 
              nn4693, nn4692, nn4691, nn4690, nn4689, nn4688, nn4687, nn4686, 
              nn4685} ), 
        .SUM( {\inputctrl1_u109_XORCI_16|SUM_net , 
              \inputctrl1_u109_XORCI_15|SUM_net , \inputctrl1_u109_XORCI_14|SUM_net , 
              \inputctrl1_u109_XORCI_13|SUM_net , \inputctrl1_u109_XORCI_12|SUM_net , 
              \inputctrl1_u109_XORCI_11|SUM_net , \inputctrl1_u109_XORCI_10|SUM_net , 
              \inputctrl1_u109_XORCI_9|SUM_net , \inputctrl1_u109_XORCI_8|SUM_net , 
              \inputctrl1_u109_XORCI_7|SUM_net , \inputctrl1_u109_XORCI_6|SUM_net , 
              \inputctrl1_u109_XORCI_5|SUM_net , \inputctrl1_u109_XORCI_4|SUM_net , 
              \inputctrl1_u109_XORCI_3|SUM_net , \inputctrl1_u109_XORCI_2|SUM_net , 
              \inputctrl1_u109_XORCI_1|SUM_net , \inputctrl1_u109_XORCI_0|SUM_net } )
      );
    CS_REGA_PRIM cal1_HS__reg ( .CLK( clkb ), .D( nn1328 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( HS_1863_net ) );
      defparam cal1_HS__reg.INIT = 0;
      defparam cal1_HS__reg.PLACE_LOCATION = "NONE";
      defparam cal1_HS__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_VSNormal__reg ( .CLK( clkb ), .D( nn1330 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \cal1_VSNormal__reg|Q_net  ) );
      defparam cal1_VSNormal__reg.INIT = 0;
      defparam cal1_VSNormal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_VSNormal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_enforceJmp__reg ( .CLK( clkb ), .D( a_acc_en_cal1_u134_mac ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \cal1_enforceJmp__reg|Q_net  ) );
      defparam cal1_enforceJmp__reg.INIT = 0;
      defparam cal1_enforceJmp__reg.PLACE_LOCATION = "NONE";
      defparam cal1_enforceJmp__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_jmp1Normal__reg ( .CLK( clkb ), .D( nn2710 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \cal1_jmp1Normal__reg|Q_net  ) );
      defparam cal1_jmp1Normal__reg.INIT = 0;
      defparam cal1_jmp1Normal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_jmp1Normal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_jmp2Normal__reg ( .CLK( clkb ), .D( nn2711 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \cal1_jmp2Normal__reg|Q_net  ) );
      defparam cal1_jmp2Normal__reg.INIT = 0;
      defparam cal1_jmp2Normal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_jmp2Normal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[0]  ( .CLK( clkb ), .D( nn4091 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[0]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[0] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[10]  ( .CLK( clkb ), .D( nn4118 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[10]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[10] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[1]  ( .CLK( clkb ), .D( nn4119 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[1]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[1] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[2]  ( .CLK( clkb ), .D( nn4120 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[2]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[2] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[3]  ( .CLK( clkb ), .D( nn4121 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[3]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[3] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[4]  ( .CLK( clkb ), .D( nn4122 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[4]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[4] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[5]  ( .CLK( clkb ), .D( nn4123 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[5]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[5] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[6]  ( .CLK( clkb ), .D( nn4124 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[6]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[6] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[7]  ( .CLK( clkb ), .D( nn4125 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[7]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[7] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[8]  ( .CLK( clkb ), .D( nn4126 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[8]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[8] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[9]  ( .CLK( clkb ), .D( nn4127 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4093 ), .Q( \cal1_ramRdAddr__reg[9]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[9] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[0]  ( .CLK( clkb ), .D( \cal1_u__reg[0]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[0]|Q_net  ) );
      defparam \cal1_uPreF__reg[0] .INIT = 0;
      defparam \cal1_uPreF__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[1]  ( .CLK( clkb ), .D( \cal1_u__reg[1]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[1]|Q_net  ) );
      defparam \cal1_uPreF__reg[1] .INIT = 0;
      defparam \cal1_uPreF__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[2]  ( .CLK( clkb ), .D( \cal1_u__reg[2]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[2]|Q_net  ) );
      defparam \cal1_uPreF__reg[2] .INIT = 0;
      defparam \cal1_uPreF__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[3]  ( .CLK( clkb ), .D( \cal1_u__reg[3]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[3]|Q_net  ) );
      defparam \cal1_uPreF__reg[3] .INIT = 0;
      defparam \cal1_uPreF__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[4]  ( .CLK( clkb ), .D( \cal1_u__reg[4]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[4]|Q_net  ) );
      defparam \cal1_uPreF__reg[4] .INIT = 0;
      defparam \cal1_uPreF__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[5]  ( .CLK( clkb ), .D( \cal1_u__reg[5]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_uPreF__reg[5]|Q_net  ) );
      defparam \cal1_uPreF__reg[5] .INIT = 0;
      defparam \cal1_uPreF__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[0]  ( .CLK( clkb ), .D( nn4129 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[0]|Q_net  ) );
      defparam \cal1_u__reg[0] .INIT = 0;
      defparam \cal1_u__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[10]  ( .CLK( clkb ), .D( nn4130 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[10]|Q_net  ) );
      defparam \cal1_u__reg[10] .INIT = 0;
      defparam \cal1_u__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[11]  ( .CLK( clkb ), .D( nn4131 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[11]|Q_net  ) );
      defparam \cal1_u__reg[11] .INIT = 0;
      defparam \cal1_u__reg[11] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[12]  ( .CLK( clkb ), .D( nn4132 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[12]|Q_net  ) );
      defparam \cal1_u__reg[12] .INIT = 0;
      defparam \cal1_u__reg[12] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[13]  ( .CLK( clkb ), .D( nn4133 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[13]|Q_net  ) );
      defparam \cal1_u__reg[13] .INIT = 0;
      defparam \cal1_u__reg[13] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[14]  ( .CLK( clkb ), .D( nn4134 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[14]|Q_net  ) );
      defparam \cal1_u__reg[14] .INIT = 0;
      defparam \cal1_u__reg[14] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[15]  ( .CLK( clkb ), .D( nn4135 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[15]|Q_net  ) );
      defparam \cal1_u__reg[15] .INIT = 0;
      defparam \cal1_u__reg[15] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[16]  ( .CLK( clkb ), .D( nn4136 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[16]|Q_net  ) );
      defparam \cal1_u__reg[16] .INIT = 0;
      defparam \cal1_u__reg[16] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[1]  ( .CLK( clkb ), .D( nn4137 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[1]|Q_net  ) );
      defparam \cal1_u__reg[1] .INIT = 0;
      defparam \cal1_u__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[2]  ( .CLK( clkb ), .D( nn4138 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[2]|Q_net  ) );
      defparam \cal1_u__reg[2] .INIT = 0;
      defparam \cal1_u__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[3]  ( .CLK( clkb ), .D( nn4139 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[3]|Q_net  ) );
      defparam \cal1_u__reg[3] .INIT = 0;
      defparam \cal1_u__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[4]  ( .CLK( clkb ), .D( nn4140 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[4]|Q_net  ) );
      defparam \cal1_u__reg[4] .INIT = 0;
      defparam \cal1_u__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[5]  ( .CLK( clkb ), .D( nn4141 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[5]|Q_net  ) );
      defparam \cal1_u__reg[5] .INIT = 0;
      defparam \cal1_u__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[6]  ( .CLK( clkb ), .D( nn4142 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[6]|Q_net  ) );
      defparam \cal1_u__reg[6] .INIT = 0;
      defparam \cal1_u__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[7]  ( .CLK( clkb ), .D( nn4143 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[7]|Q_net  ) );
      defparam \cal1_u__reg[7] .INIT = 0;
      defparam \cal1_u__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[8]  ( .CLK( clkb ), .D( nn4144 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[8]|Q_net  ) );
      defparam \cal1_u__reg[8] .INIT = 0;
      defparam \cal1_u__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[9]  ( .CLK( clkb ), .D( nn4145 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_u__reg[9]|Q_net  ) );
      defparam \cal1_u__reg[9] .INIT = 0;
      defparam \cal1_u__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[0]  ( .CLK( clkb ), .D( nn4147 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[0]|Q_net  ) );
      defparam \cal1_v__reg[0] .INIT = 0;
      defparam \cal1_v__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[10]  ( .CLK( clkb ), .D( nn4148 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[10]|Q_net  ) );
      defparam \cal1_v__reg[10] .INIT = 0;
      defparam \cal1_v__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[11]  ( .CLK( clkb ), .D( nn4149 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[11]|Q_net  ) );
      defparam \cal1_v__reg[11] .INIT = 0;
      defparam \cal1_v__reg[11] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[12]  ( .CLK( clkb ), .D( nn4150 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[12]|Q_net  ) );
      defparam \cal1_v__reg[12] .INIT = 0;
      defparam \cal1_v__reg[12] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[13]  ( .CLK( clkb ), .D( nn4151 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[13]|Q_net  ) );
      defparam \cal1_v__reg[13] .INIT = 0;
      defparam \cal1_v__reg[13] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[14]  ( .CLK( clkb ), .D( nn4152 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[14]|Q_net  ) );
      defparam \cal1_v__reg[14] .INIT = 0;
      defparam \cal1_v__reg[14] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[15]  ( .CLK( clkb ), .D( nn4153 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[15]|Q_net  ) );
      defparam \cal1_v__reg[15] .INIT = 0;
      defparam \cal1_v__reg[15] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[16]  ( .CLK( clkb ), .D( nn4154 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[16]|Q_net  ) );
      defparam \cal1_v__reg[16] .INIT = 0;
      defparam \cal1_v__reg[16] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[1]  ( .CLK( clkb ), .D( nn4155 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[1]|Q_net  ) );
      defparam \cal1_v__reg[1] .INIT = 0;
      defparam \cal1_v__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[2]  ( .CLK( clkb ), .D( nn4156 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[2]|Q_net  ) );
      defparam \cal1_v__reg[2] .INIT = 0;
      defparam \cal1_v__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[3]  ( .CLK( clkb ), .D( nn4157 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[3]|Q_net  ) );
      defparam \cal1_v__reg[3] .INIT = 0;
      defparam \cal1_v__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[4]  ( .CLK( clkb ), .D( nn4158 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[4]|Q_net  ) );
      defparam \cal1_v__reg[4] .INIT = 0;
      defparam \cal1_v__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[5]  ( .CLK( clkb ), .D( nn4159 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[5]|Q_net  ) );
      defparam \cal1_v__reg[5] .INIT = 0;
      defparam \cal1_v__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[6]  ( .CLK( clkb ), .D( nn4160 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[6]|Q_net  ) );
      defparam \cal1_v__reg[6] .INIT = 0;
      defparam \cal1_v__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[7]  ( .CLK( clkb ), .D( nn4161 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[7]|Q_net  ) );
      defparam \cal1_v__reg[7] .INIT = 0;
      defparam \cal1_v__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[8]  ( .CLK( clkb ), .D( nn4162 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[8]|Q_net  ) );
      defparam \cal1_v__reg[8] .INIT = 0;
      defparam \cal1_v__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[9]  ( .CLK( clkb ), .D( nn4163 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_v__reg[9]|Q_net  ) );
      defparam \cal1_v__reg[9] .INIT = 0;
      defparam \cal1_v__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[0]  ( .CLK( clkb ), .D( nn4164 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[0]|Q_net  ) );
      defparam \cal1_xAddress__reg[0] .INIT = 0;
      defparam \cal1_xAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[10]  ( .CLK( clkb ), .D( nn4189 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[10]|Q_net  ) );
      defparam \cal1_xAddress__reg[10] .INIT = 0;
      defparam \cal1_xAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[1]  ( .CLK( clkb ), .D( nn4190 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[1]|Q_net  ) );
      defparam \cal1_xAddress__reg[1] .INIT = 0;
      defparam \cal1_xAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[2]  ( .CLK( clkb ), .D( nn4191 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[2]|Q_net  ) );
      defparam \cal1_xAddress__reg[2] .INIT = 0;
      defparam \cal1_xAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[3]  ( .CLK( clkb ), .D( nn4192 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[3]|Q_net  ) );
      defparam \cal1_xAddress__reg[3] .INIT = 0;
      defparam \cal1_xAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[4]  ( .CLK( clkb ), .D( nn4193 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[4]|Q_net  ) );
      defparam \cal1_xAddress__reg[4] .INIT = 0;
      defparam \cal1_xAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[5]  ( .CLK( clkb ), .D( nn4194 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[5]|Q_net  ) );
      defparam \cal1_xAddress__reg[5] .INIT = 0;
      defparam \cal1_xAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[6]  ( .CLK( clkb ), .D( nn4195 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[6]|Q_net  ) );
      defparam \cal1_xAddress__reg[6] .INIT = 0;
      defparam \cal1_xAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[7]  ( .CLK( clkb ), .D( nn4196 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[7]|Q_net  ) );
      defparam \cal1_xAddress__reg[7] .INIT = 0;
      defparam \cal1_xAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[8]  ( .CLK( clkb ), .D( nn4197 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[8]|Q_net  ) );
      defparam \cal1_xAddress__reg[8] .INIT = 0;
      defparam \cal1_xAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[9]  ( .CLK( clkb ), .D( nn4198 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4092 ), .Q( \cal1_xAddress__reg[9]|Q_net  ) );
      defparam \cal1_xAddress__reg[9] .INIT = 0;
      defparam \cal1_xAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[0]  ( .CLK( clkb ), .D( nn4199 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[0]|Q_net  ) );
      defparam \cal1_yAddress__reg[0] .INIT = 0;
      defparam \cal1_yAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[10]  ( .CLK( clkb ), .D( nn4224 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[10]|Q_net  ) );
      defparam \cal1_yAddress__reg[10] .INIT = 0;
      defparam \cal1_yAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[1]  ( .CLK( clkb ), .D( nn4225 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[1]|Q_net  ) );
      defparam \cal1_yAddress__reg[1] .INIT = 0;
      defparam \cal1_yAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[2]  ( .CLK( clkb ), .D( nn4226 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[2]|Q_net  ) );
      defparam \cal1_yAddress__reg[2] .INIT = 0;
      defparam \cal1_yAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[3]  ( .CLK( clkb ), .D( nn4227 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[3]|Q_net  ) );
      defparam \cal1_yAddress__reg[3] .INIT = 0;
      defparam \cal1_yAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[4]  ( .CLK( clkb ), .D( nn4228 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[4]|Q_net  ) );
      defparam \cal1_yAddress__reg[4] .INIT = 0;
      defparam \cal1_yAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[5]  ( .CLK( clkb ), .D( nn4229 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[5]|Q_net  ) );
      defparam \cal1_yAddress__reg[5] .INIT = 0;
      defparam \cal1_yAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[6]  ( .CLK( clkb ), .D( nn4230 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[6]|Q_net  ) );
      defparam \cal1_yAddress__reg[6] .INIT = 0;
      defparam \cal1_yAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[7]  ( .CLK( clkb ), .D( nn4231 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[7]|Q_net  ) );
      defparam \cal1_yAddress__reg[7] .INIT = 0;
      defparam \cal1_yAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[8]  ( .CLK( clkb ), .D( nn4232 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[8]|Q_net  ) );
      defparam \cal1_yAddress__reg[8] .INIT = 0;
      defparam \cal1_yAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[9]  ( .CLK( clkb ), .D( nn4233 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn1329 ), .Q( \cal1_yAddress__reg[9]|Q_net  ) );
      defparam \cal1_yAddress__reg[9] .INIT = 0;
      defparam \cal1_yAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[0]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[0] .INIT = 0;
      defparam \coefcal1_frameRate__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[1]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[1] .INIT = 0;
      defparam \coefcal1_frameRate__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[2]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[2]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[2] .INIT = 0;
      defparam \coefcal1_frameRate__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[3]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[3] .INIT = 0;
      defparam \coefcal1_frameRate__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[4]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[4] .INIT = 0;
      defparam \coefcal1_frameRate__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[5]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[5]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[5] .INIT = 0;
      defparam \coefcal1_frameRate__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[6]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[6]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[6] .INIT = 0;
      defparam \coefcal1_frameRate__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[7]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[7]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[7] .INIT = 0;
      defparam \coefcal1_frameRate__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[8]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_frameRate__reg[8]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[8] .INIT = 0;
      defparam \coefcal1_frameRate__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM coefcal1_inEn__reg ( .CLK( clka ), .D( nn4234 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_inEn__reg|Q_net  ) );
      defparam coefcal1_inEn__reg.INIT = 0;
      defparam coefcal1_inEn__reg.PLACE_LOCATION = "NONE";
      defparam coefcal1_inEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM coefcal1_work__reg ( .CLK( clka ), .D( nn4336 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_work__reg|Q_net  ) );
      defparam coefcal1_work__reg.INIT = 0;
      defparam coefcal1_work__reg.PLACE_LOCATION = "NONE";
      defparam coefcal1_work__reg.PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[0]|Q_net  ) );
      defparam \coefcal1_working__reg[0] .INIT = 0;
      defparam \coefcal1_working__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[10]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[10]|Q_net  ) );
      defparam \coefcal1_working__reg[10] .INIT = 0;
      defparam \coefcal1_working__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[11]|Q_net  ) );
      defparam \coefcal1_working__reg[11] .INIT = 0;
      defparam \coefcal1_working__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[12]|Q_net  ) );
      defparam \coefcal1_working__reg[12] .INIT = 0;
      defparam \coefcal1_working__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[13]|Q_net  ) );
      defparam \coefcal1_working__reg[13] .INIT = 0;
      defparam \coefcal1_working__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[14]|Q_net  ) );
      defparam \coefcal1_working__reg[14] .INIT = 0;
      defparam \coefcal1_working__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[15]|Q_net  ) );
      defparam \coefcal1_working__reg[15] .INIT = 0;
      defparam \coefcal1_working__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[16]|Q_net  ) );
      defparam \coefcal1_working__reg[16] .INIT = 0;
      defparam \coefcal1_working__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[17]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[17]|Q_net  ) );
      defparam \coefcal1_working__reg[17] .INIT = 0;
      defparam \coefcal1_working__reg[17] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[17] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[18]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[18]|Q_net  ) );
      defparam \coefcal1_working__reg[18] .INIT = 0;
      defparam \coefcal1_working__reg[18] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[18] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[19]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[19]|Q_net  ) );
      defparam \coefcal1_working__reg[19] .INIT = 0;
      defparam \coefcal1_working__reg[19] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[19] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[1]|Q_net  ) );
      defparam \coefcal1_working__reg[1] .INIT = 0;
      defparam \coefcal1_working__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[20]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[20]|Q_net  ) );
      defparam \coefcal1_working__reg[20] .INIT = 0;
      defparam \coefcal1_working__reg[20] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[20] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[21]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[21]|Q_net  ) );
      defparam \coefcal1_working__reg[21] .INIT = 0;
      defparam \coefcal1_working__reg[21] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[21] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[22]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[22]|Q_net  ) );
      defparam \coefcal1_working__reg[22] .INIT = 0;
      defparam \coefcal1_working__reg[22] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[22] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[23]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[23]|Q_net  ) );
      defparam \coefcal1_working__reg[23] .INIT = 0;
      defparam \coefcal1_working__reg[23] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[23] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[24]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[24]|Q_net  ) );
      defparam \coefcal1_working__reg[24] .INIT = 0;
      defparam \coefcal1_working__reg[24] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[24] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[25]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[25]|Q_net  ) );
      defparam \coefcal1_working__reg[25] .INIT = 0;
      defparam \coefcal1_working__reg[25] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[25] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[26]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[26]|Q_net  ) );
      defparam \coefcal1_working__reg[26] .INIT = 0;
      defparam \coefcal1_working__reg[26] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[26] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[27]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[27]|Q_net  ) );
      defparam \coefcal1_working__reg[27] .INIT = 0;
      defparam \coefcal1_working__reg[27] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[27] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[28]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[28]|Q_net  ) );
      defparam \coefcal1_working__reg[28] .INIT = 0;
      defparam \coefcal1_working__reg[28] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[28] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[29]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[29]|Q_net  ) );
      defparam \coefcal1_working__reg[29] .INIT = 0;
      defparam \coefcal1_working__reg[29] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[29] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[2]|Q_net  ) );
      defparam \coefcal1_working__reg[2] .INIT = 0;
      defparam \coefcal1_working__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[30]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[30]|Q_net  ) );
      defparam \coefcal1_working__reg[30] .INIT = 0;
      defparam \coefcal1_working__reg[30] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[30] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[31]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[31]|Q_net  ) );
      defparam \coefcal1_working__reg[31] .INIT = 0;
      defparam \coefcal1_working__reg[31] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[31] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[32]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[32]|Q_net  ) );
      defparam \coefcal1_working__reg[32] .INIT = 0;
      defparam \coefcal1_working__reg[32] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[32] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[3]|Q_net  ) );
      defparam \coefcal1_working__reg[3] .INIT = 0;
      defparam \coefcal1_working__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[4]|Q_net  ) );
      defparam \coefcal1_working__reg[4] .INIT = 0;
      defparam \coefcal1_working__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[5]|Q_net  ) );
      defparam \coefcal1_working__reg[5] .INIT = 0;
      defparam \coefcal1_working__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[6]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[6]|Q_net  ) );
      defparam \coefcal1_working__reg[6] .INIT = 0;
      defparam \coefcal1_working__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[7]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[7]|Q_net  ) );
      defparam \coefcal1_working__reg[7] .INIT = 0;
      defparam \coefcal1_working__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[8]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[8]|Q_net  ) );
      defparam \coefcal1_working__reg[8] .INIT = 0;
      defparam \coefcal1_working__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[9]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_working__reg[9]|Q_net  ) );
      defparam \coefcal1_working__reg[9] .INIT = 0;
      defparam \coefcal1_working__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[0]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[0] .INIT = 0;
      defparam \coefcal1_xDividend__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[10]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_4|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[10]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[10] .INIT = 0;
      defparam \coefcal1_xDividend__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[11]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_5|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[11]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[11] .INIT = 0;
      defparam \coefcal1_xDividend__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[12]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_6|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[12]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[12] .INIT = 0;
      defparam \coefcal1_xDividend__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[13]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_7|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[13]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[13] .INIT = 0;
      defparam \coefcal1_xDividend__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[14]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_8|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[14]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[14] .INIT = 0;
      defparam \coefcal1_xDividend__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[15]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_9|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[15]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[15] .INIT = 0;
      defparam \coefcal1_xDividend__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[16]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[16]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[16] .INIT = 0;
      defparam \coefcal1_xDividend__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[1]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[1] .INIT = 0;
      defparam \coefcal1_xDividend__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[2]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[2] .INIT = 0;
      defparam \coefcal1_xDividend__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[3]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[3] .INIT = 0;
      defparam \coefcal1_xDividend__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[4]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[4] .INIT = 0;
      defparam \coefcal1_xDividend__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[5]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[5] .INIT = 0;
      defparam \coefcal1_xDividend__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[6]  ( .CLK( clka ), .D( nn4361 ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[6]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[6] .INIT = 0;
      defparam \coefcal1_xDividend__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[7]  ( .CLK( clka ), .D( nn4362 ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[7]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[7] .INIT = 0;
      defparam \coefcal1_xDividend__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[8]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_2|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[8]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[8] .INIT = 0;
      defparam \coefcal1_xDividend__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[9]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_3|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDividend__reg[9]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[9] .INIT = 0;
      defparam \coefcal1_xDividend__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[0]  ( .CLK( clka ), .D( outXRes[0] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[0]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[0] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[10]  ( .CLK( clka ), .D( outXRes[10] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[10]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[10] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[11]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[11] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[12]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[12] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[13]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[13] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[14]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[14] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[15]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[15] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[16]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[16] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[1]  ( .CLK( clka ), .D( outXRes[1] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[1]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[1] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[2]  ( .CLK( clka ), .D( outXRes[2] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[2]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[2] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[3]  ( .CLK( clka ), .D( outXRes[3] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[3]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[3] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[4]  ( .CLK( clka ), .D( outXRes[4] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[4]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[4] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[5]  ( .CLK( clka ), .D( outXRes[5] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[5]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[5] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[6]  ( .CLK( clka ), .D( outXRes[6] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[6]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[6] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[7]  ( .CLK( clka ), .D( outXRes[7] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[7]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[7] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[8]  ( .CLK( clka ), .D( outXRes[8] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[8]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[8] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[9]  ( .CLK( clka ), .D( outXRes[9] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_xDivisor__reg[9]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[9] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[0]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[0] .INIT = 0;
      defparam \coefcal1_yDividend__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[10]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_4|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[10]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[10] .INIT = 0;
      defparam \coefcal1_yDividend__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[11]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_5|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[11]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[11] .INIT = 0;
      defparam \coefcal1_yDividend__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[12]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_6|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[12]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[12] .INIT = 0;
      defparam \coefcal1_yDividend__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[13]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_7|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[13]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[13] .INIT = 0;
      defparam \coefcal1_yDividend__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[14]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_8|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[14]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[14] .INIT = 0;
      defparam \coefcal1_yDividend__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[15]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_9|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[15]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[15] .INIT = 0;
      defparam \coefcal1_yDividend__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[16]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[16]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[16] .INIT = 0;
      defparam \coefcal1_yDividend__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[1]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[1] .INIT = 0;
      defparam \coefcal1_yDividend__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[2]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[2] .INIT = 0;
      defparam \coefcal1_yDividend__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[3]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[3] .INIT = 0;
      defparam \coefcal1_yDividend__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[4]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[4] .INIT = 0;
      defparam \coefcal1_yDividend__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[5]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[5] .INIT = 0;
      defparam \coefcal1_yDividend__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[6]  ( .CLK( clka ), .D( nn4413 ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[6]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[6] .INIT = 0;
      defparam \coefcal1_yDividend__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[7]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_1|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[7]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[7] .INIT = 0;
      defparam \coefcal1_yDividend__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[8]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_2|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[8]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[8] .INIT = 0;
      defparam \coefcal1_yDividend__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[9]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_3|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDividend__reg[9]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[9] .INIT = 0;
      defparam \coefcal1_yDividend__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[0]  ( .CLK( clka ), .D( outYRes[0] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[0]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[0] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[10]  ( .CLK( clka ), .D( outYRes[10] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[10]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[10] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[11]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[11] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[12]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[12] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[13]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[13] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[14]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[14] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[15]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[15] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u134_mac ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[16]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[16] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[1]  ( .CLK( clka ), .D( outYRes[1] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[1]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[1] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[2]  ( .CLK( clka ), .D( outYRes[2] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[2]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[2] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[3]  ( .CLK( clka ), .D( outYRes[3] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[3]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[3] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[4]  ( .CLK( clka ), .D( outYRes[4] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[4]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[4] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[5]  ( .CLK( clka ), .D( outYRes[5] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[5]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[5] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[6]  ( .CLK( clka ), .D( outYRes[6] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[6]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[6] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[7]  ( .CLK( clka ), .D( outYRes[7] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[7]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[7] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[8]  ( .CLK( clka ), .D( outYRes[8] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[8]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[8] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[9]  ( .CLK( clka ), .D( outYRes[9] ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \coefcal1_yDivisor__reg[9]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[9] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_0_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_0_u_emb18k_0  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_0_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_0_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1_u_emb18k_0  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_1_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_1_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1_u_emb18k_0  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_3_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u134_mac ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \fifo1_ram_inst_3_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[0]  ( .CLK( clka ), .D( nn4414 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[0]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[0] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[10]  ( .CLK( clka ), .D( nn4537 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[10]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[10] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[11]  ( .CLK( clka ), .D( nn4538 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[11]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[11] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[12]  ( .CLK( clka ), .D( nn4539 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[12]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[12] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[13]  ( .CLK( clka ), .D( nn4540 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[13]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[13] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[14]  ( .CLK( clka ), .D( nn4541 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[14]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[14] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[15]  ( .CLK( clka ), .D( nn4542 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[15]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[15] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[1]  ( .CLK( clka ), .D( nn4543 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[1]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[1] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[2]  ( .CLK( clka ), .D( nn4544 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[2]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[2] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[3]  ( .CLK( clka ), .D( nn4545 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[3]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[3] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[4]  ( .CLK( clka ), .D( nn4546 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[4]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[4] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[5]  ( .CLK( clka ), .D( nn4547 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[5]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[5] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[6]  ( .CLK( clka ), .D( nn4548 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[6]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[6] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[7]  ( .CLK( clka ), .D( nn4549 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[7]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[7] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[8]  ( .CLK( clka ), .D( nn4550 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[8]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[8] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[9]  ( .CLK( clka ), .D( nn4551 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_dataOut__reg[9]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[9] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_jmp__reg ( .CLK( clka ), .D( nn4552 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4536 ), .Q( \inputctrl1_jmp__reg|Q_net  ) );
      defparam inputctrl1_jmp__reg.INIT = 0;
      defparam inputctrl1_jmp__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_jmp__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[0]  ( .CLK( clka ), .D( nn4553 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[0]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[0] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[10]  ( .CLK( clka ), .D( nn4578 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[10]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[10] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[1]  ( .CLK( clka ), .D( nn4579 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[1]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[1] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[2]  ( .CLK( clka ), .D( nn4580 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[2]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[2] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[3]  ( .CLK( clka ), .D( nn4581 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[3]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[3] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[4]  ( .CLK( clka ), .D( nn4582 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[4]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[4] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[5]  ( .CLK( clka ), .D( nn4583 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[5]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[5] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[6]  ( .CLK( clka ), .D( nn4584 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[6]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[6] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[7]  ( .CLK( clka ), .D( nn4585 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[7]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[7] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[8]  ( .CLK( clka ), .D( nn4586 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[8]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[8] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[9]  ( .CLK( clka ), .D( nn4587 ), .RST( a_acc_en_cal1_u134_mac ), .SET( rst ), .CE( nn4536 ), .Q( \inputctrl1_ramWrtAddr__reg[9]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[9] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_ramWrtEn__reg ( .CLK( clka ), .D( nn4588 ), .RST( rst ), .SET( a_acc_en_cal1_u134_mac ), .CE( a_dinxy_cen_cal1_u134_mac ), .Q( \inputctrl1_ramWrtEn__reg|Q_net  ) );
      defparam inputctrl1_ramWrtEn__reg.INIT = 0;
      defparam inputctrl1_ramWrtEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_ramWrtEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[0]  ( .CLK( clka ), .D( nn4589 ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[0]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[0] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_10|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[10]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[10] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_1|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[1]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[1] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_2|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[2]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[2] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_3|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[3]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[3] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_4|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[4]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[4] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_5|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[5]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[5] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_6|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[6]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[6] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_7|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[7]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[7] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_8|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[8]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[8] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_9|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xAddress__reg[9]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[9] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[0]  ( .CLK( clka ), .D( nn4617 ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[0]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[0] .INIT = 0;
      defparam \inputctrl1_xCal__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_10|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[10]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[10] .INIT = 0;
      defparam \inputctrl1_xCal__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[11]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_11|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[11]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[11] .INIT = 0;
      defparam \inputctrl1_xCal__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[12]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_12|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[12]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[12] .INIT = 0;
      defparam \inputctrl1_xCal__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[13]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_13|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[13]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[13] .INIT = 0;
      defparam \inputctrl1_xCal__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[14]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_14|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[14]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[14] .INIT = 0;
      defparam \inputctrl1_xCal__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[15]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_15|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[15]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[15] .INIT = 0;
      defparam \inputctrl1_xCal__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[16]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_16|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[16]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[16] .INIT = 0;
      defparam \inputctrl1_xCal__reg[16] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_1|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[1]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[1] .INIT = 0;
      defparam \inputctrl1_xCal__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_2|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[2]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[2] .INIT = 0;
      defparam \inputctrl1_xCal__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_3|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[3]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[3] .INIT = 0;
      defparam \inputctrl1_xCal__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_4|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[4]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[4] .INIT = 0;
      defparam \inputctrl1_xCal__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_5|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[5]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[5] .INIT = 0;
      defparam \inputctrl1_xCal__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_6|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[6]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[6] .INIT = 0;
      defparam \inputctrl1_xCal__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_7|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[7]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[7] .INIT = 0;
      defparam \inputctrl1_xCal__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_8|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[8]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[8] .INIT = 0;
      defparam \inputctrl1_xCal__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_9|SUM_net  ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4618 ), .Q( \inputctrl1_xCal__reg[9]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[9] .INIT = 0;
      defparam \inputctrl1_xCal__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_xPreEn__reg ( .CLK( clka ), .D( nn4455 ), .RST( nn4590 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4591 ), .Q( \inputctrl1_xPreEn__reg|Q_net  ) );
      defparam inputctrl1_xPreEn__reg.INIT = 0;
      defparam inputctrl1_xPreEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_xPreEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[0]  ( .CLK( clka ), .D( nn4655 ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[0]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[0] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_10|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[10]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[10] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_1|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[1]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[1] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_2|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[2]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[2] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_3|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[3]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[3] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_4|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[4]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[4] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_5|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[5]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[5] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_6|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[6]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[6] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_7|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[7]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[7] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_8|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[8]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[8] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_9|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[9]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[9] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[0]  ( .CLK( clka ), .D( nn4683 ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[0]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[0] .INIT = 0;
      defparam \inputctrl1_yCal__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_10|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[10]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[10] .INIT = 0;
      defparam \inputctrl1_yCal__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[11]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_11|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[11]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[11] .INIT = 0;
      defparam \inputctrl1_yCal__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[12]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_12|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[12]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[12] .INIT = 0;
      defparam \inputctrl1_yCal__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[13]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_13|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[13]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[13] .INIT = 0;
      defparam \inputctrl1_yCal__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[14]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_14|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[14]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[14] .INIT = 0;
      defparam \inputctrl1_yCal__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[15]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_15|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[15]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[15] .INIT = 0;
      defparam \inputctrl1_yCal__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[16]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_16|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[16]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[16] .INIT = 0;
      defparam \inputctrl1_yCal__reg[16] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_1|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[1]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[1] .INIT = 0;
      defparam \inputctrl1_yCal__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_2|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[2]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[2] .INIT = 0;
      defparam \inputctrl1_yCal__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_3|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[3]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[3] .INIT = 0;
      defparam \inputctrl1_yCal__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_4|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[4]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[4] .INIT = 0;
      defparam \inputctrl1_yCal__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_5|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[5]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[5] .INIT = 0;
      defparam \inputctrl1_yCal__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_6|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[6]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[6] .INIT = 0;
      defparam \inputctrl1_yCal__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_7|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[7]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[7] .INIT = 0;
      defparam \inputctrl1_yCal__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_8|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[8]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[8] .INIT = 0;
      defparam \inputctrl1_yCal__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_9|SUM_net  ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( nn4684 ), .Q( \inputctrl1_yCal__reg[9]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[9] .INIT = 0;
      defparam \inputctrl1_yCal__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_yPreEn__reg ( .CLK( clka ), .D( nn4421 ), .RST( nn4656 ), .SET( a_acc_en_cal1_u134_mac ), .CE( iHsyn ), .Q( \inputctrl1_yPreEn__reg|Q_net  ) );
      defparam inputctrl1_yPreEn__reg.INIT = 0;
      defparam inputctrl1_yPreEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_yPreEn__reg.PCK_LOCATION = "NONE";

endmodule


