module scaler_ipc_adder_10(CA, CI, CO, DX, SUM);
  input [9:0] CA;
  input CI;
  output CO;
  input [9:0] DX;
  output [9:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(CO), 
        .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_11(CA, CI, CO, DX, SUM);
  input [10:0] CA;
  input CI;
  output CO;
  input [10:0] DX;
  output [10:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(CO), 
        .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_12(CA, CI, CO, DX, SUM);
  input [11:0] CA;
  input CI;
  output CO;
  input [11:0] DX;
  output [11:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(CO), 
        .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_14(CA, CI, CO, DX, SUM);
  input [13:0] CA;
  input CI;
  output CO;
  input [13:0] DX;
  output [13:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(CO), 
        .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_17(CA, CI, CO, DX, SUM);
  input [16:0] CA;
  input CI;
  output CO;
  input [16:0] DX;
  output [16:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(CO), 
        .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_18(CA, CI, CO, DX, SUM);
  input [17:0] CA;
  input CI;
  output CO;
  input [17:0] DX;
  output [17:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_16|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(
        \MUXCO_16|COUT_net ), .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_17 ( .AIN(CA[17]), .CIN(\MUXCO_16|COUT_net ), .COUT(CO), 
        .CSEL(DX[17]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_17 ( .CIN(\MUXCO_16|COUT_net ), .DIN(DX[17]), .SUM(
        SUM[17]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_34(CA, CI, CO, DX, SUM);
  input [33:0] CA;
  input CI;
  output CO;
  input [33:0] DX;
  output [33:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_10|COUT_net ;
    wire \MUXCO_11|COUT_net ;
    wire \MUXCO_12|COUT_net ;
    wire \MUXCO_13|COUT_net ;
    wire \MUXCO_14|COUT_net ;
    wire \MUXCO_15|COUT_net ;
    wire \MUXCO_16|COUT_net ;
    wire \MUXCO_17|COUT_net ;
    wire \MUXCO_18|COUT_net ;
    wire \MUXCO_19|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_20|COUT_net ;
    wire \MUXCO_21|COUT_net ;
    wire \MUXCO_22|COUT_net ;
    wire \MUXCO_23|COUT_net ;
    wire \MUXCO_24|COUT_net ;
    wire \MUXCO_25|COUT_net ;
    wire \MUXCO_26|COUT_net ;
    wire \MUXCO_27|COUT_net ;
    wire \MUXCO_28|COUT_net ;
    wire \MUXCO_29|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_30|COUT_net ;
    wire \MUXCO_31|COUT_net ;
    wire \MUXCO_32|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;
    wire \MUXCO_8|COUT_net ;
    wire \MUXCO_9|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_10 ( .AIN(CA[10]), .CIN(\MUXCO_9|COUT_net ), .COUT(
        \MUXCO_10|COUT_net ), .CSEL(DX[10]) );
    CS_MUXCO_PRIM MUXCO_11 ( .AIN(CA[11]), .CIN(\MUXCO_10|COUT_net ), .COUT(
        \MUXCO_11|COUT_net ), .CSEL(DX[11]) );
    CS_MUXCO_PRIM MUXCO_12 ( .AIN(CA[12]), .CIN(\MUXCO_11|COUT_net ), .COUT(
        \MUXCO_12|COUT_net ), .CSEL(DX[12]) );
    CS_MUXCO_PRIM MUXCO_13 ( .AIN(CA[13]), .CIN(\MUXCO_12|COUT_net ), .COUT(
        \MUXCO_13|COUT_net ), .CSEL(DX[13]) );
    CS_MUXCO_PRIM MUXCO_14 ( .AIN(CA[14]), .CIN(\MUXCO_13|COUT_net ), .COUT(
        \MUXCO_14|COUT_net ), .CSEL(DX[14]) );
    CS_MUXCO_PRIM MUXCO_15 ( .AIN(CA[15]), .CIN(\MUXCO_14|COUT_net ), .COUT(
        \MUXCO_15|COUT_net ), .CSEL(DX[15]) );
    CS_MUXCO_PRIM MUXCO_16 ( .AIN(CA[16]), .CIN(\MUXCO_15|COUT_net ), .COUT(
        \MUXCO_16|COUT_net ), .CSEL(DX[16]) );
    CS_MUXCO_PRIM MUXCO_17 ( .AIN(CA[17]), .CIN(\MUXCO_16|COUT_net ), .COUT(
        \MUXCO_17|COUT_net ), .CSEL(DX[17]) );
    CS_MUXCO_PRIM MUXCO_18 ( .AIN(CA[18]), .CIN(\MUXCO_17|COUT_net ), .COUT(
        \MUXCO_18|COUT_net ), .CSEL(DX[18]) );
    CS_MUXCO_PRIM MUXCO_19 ( .AIN(CA[19]), .CIN(\MUXCO_18|COUT_net ), .COUT(
        \MUXCO_19|COUT_net ), .CSEL(DX[19]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_20 ( .AIN(CA[20]), .CIN(\MUXCO_19|COUT_net ), .COUT(
        \MUXCO_20|COUT_net ), .CSEL(DX[20]) );
    CS_MUXCO_PRIM MUXCO_21 ( .AIN(CA[21]), .CIN(\MUXCO_20|COUT_net ), .COUT(
        \MUXCO_21|COUT_net ), .CSEL(DX[21]) );
    CS_MUXCO_PRIM MUXCO_22 ( .AIN(CA[22]), .CIN(\MUXCO_21|COUT_net ), .COUT(
        \MUXCO_22|COUT_net ), .CSEL(DX[22]) );
    CS_MUXCO_PRIM MUXCO_23 ( .AIN(CA[23]), .CIN(\MUXCO_22|COUT_net ), .COUT(
        \MUXCO_23|COUT_net ), .CSEL(DX[23]) );
    CS_MUXCO_PRIM MUXCO_24 ( .AIN(CA[24]), .CIN(\MUXCO_23|COUT_net ), .COUT(
        \MUXCO_24|COUT_net ), .CSEL(DX[24]) );
    CS_MUXCO_PRIM MUXCO_25 ( .AIN(CA[25]), .CIN(\MUXCO_24|COUT_net ), .COUT(
        \MUXCO_25|COUT_net ), .CSEL(DX[25]) );
    CS_MUXCO_PRIM MUXCO_26 ( .AIN(CA[26]), .CIN(\MUXCO_25|COUT_net ), .COUT(
        \MUXCO_26|COUT_net ), .CSEL(DX[26]) );
    CS_MUXCO_PRIM MUXCO_27 ( .AIN(CA[27]), .CIN(\MUXCO_26|COUT_net ), .COUT(
        \MUXCO_27|COUT_net ), .CSEL(DX[27]) );
    CS_MUXCO_PRIM MUXCO_28 ( .AIN(CA[28]), .CIN(\MUXCO_27|COUT_net ), .COUT(
        \MUXCO_28|COUT_net ), .CSEL(DX[28]) );
    CS_MUXCO_PRIM MUXCO_29 ( .AIN(CA[29]), .CIN(\MUXCO_28|COUT_net ), .COUT(
        \MUXCO_29|COUT_net ), .CSEL(DX[29]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_30 ( .AIN(CA[30]), .CIN(\MUXCO_29|COUT_net ), .COUT(
        \MUXCO_30|COUT_net ), .CSEL(DX[30]) );
    CS_MUXCO_PRIM MUXCO_31 ( .AIN(CA[31]), .CIN(\MUXCO_30|COUT_net ), .COUT(
        \MUXCO_31|COUT_net ), .CSEL(DX[31]) );
    CS_MUXCO_PRIM MUXCO_32 ( .AIN(CA[32]), .CIN(\MUXCO_31|COUT_net ), .COUT(
        \MUXCO_32|COUT_net ), .CSEL(DX[32]) );
    CS_MUXCO_PRIM MUXCO_33 ( .AIN(CA[33]), .CIN(\MUXCO_32|COUT_net ), .COUT(CO), 
        .CSEL(DX[33]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(
        \MUXCO_8|COUT_net ), .CSEL(DX[8]) );
    CS_MUXCO_PRIM MUXCO_9 ( .AIN(CA[9]), .CIN(\MUXCO_8|COUT_net ), .COUT(
        \MUXCO_9|COUT_net ), .CSEL(DX[9]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_10 ( .CIN(\MUXCO_9|COUT_net ), .DIN(DX[10]), .SUM(
        SUM[10]) );
    CS_XORCI_PRIM XORCI_11 ( .CIN(\MUXCO_10|COUT_net ), .DIN(DX[11]), .SUM(
        SUM[11]) );
    CS_XORCI_PRIM XORCI_12 ( .CIN(\MUXCO_11|COUT_net ), .DIN(DX[12]), .SUM(
        SUM[12]) );
    CS_XORCI_PRIM XORCI_13 ( .CIN(\MUXCO_12|COUT_net ), .DIN(DX[13]), .SUM(
        SUM[13]) );
    CS_XORCI_PRIM XORCI_14 ( .CIN(\MUXCO_13|COUT_net ), .DIN(DX[14]), .SUM(
        SUM[14]) );
    CS_XORCI_PRIM XORCI_15 ( .CIN(\MUXCO_14|COUT_net ), .DIN(DX[15]), .SUM(
        SUM[15]) );
    CS_XORCI_PRIM XORCI_16 ( .CIN(\MUXCO_15|COUT_net ), .DIN(DX[16]), .SUM(
        SUM[16]) );
    CS_XORCI_PRIM XORCI_17 ( .CIN(\MUXCO_16|COUT_net ), .DIN(DX[17]), .SUM(
        SUM[17]) );
    CS_XORCI_PRIM XORCI_18 ( .CIN(\MUXCO_17|COUT_net ), .DIN(DX[18]), .SUM(
        SUM[18]) );
    CS_XORCI_PRIM XORCI_19 ( .CIN(\MUXCO_18|COUT_net ), .DIN(DX[19]), .SUM(
        SUM[19]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_20 ( .CIN(\MUXCO_19|COUT_net ), .DIN(DX[20]), .SUM(
        SUM[20]) );
    CS_XORCI_PRIM XORCI_21 ( .CIN(\MUXCO_20|COUT_net ), .DIN(DX[21]), .SUM(
        SUM[21]) );
    CS_XORCI_PRIM XORCI_22 ( .CIN(\MUXCO_21|COUT_net ), .DIN(DX[22]), .SUM(
        SUM[22]) );
    CS_XORCI_PRIM XORCI_23 ( .CIN(\MUXCO_22|COUT_net ), .DIN(DX[23]), .SUM(
        SUM[23]) );
    CS_XORCI_PRIM XORCI_24 ( .CIN(\MUXCO_23|COUT_net ), .DIN(DX[24]), .SUM(
        SUM[24]) );
    CS_XORCI_PRIM XORCI_25 ( .CIN(\MUXCO_24|COUT_net ), .DIN(DX[25]), .SUM(
        SUM[25]) );
    CS_XORCI_PRIM XORCI_26 ( .CIN(\MUXCO_25|COUT_net ), .DIN(DX[26]), .SUM(
        SUM[26]) );
    CS_XORCI_PRIM XORCI_27 ( .CIN(\MUXCO_26|COUT_net ), .DIN(DX[27]), .SUM(
        SUM[27]) );
    CS_XORCI_PRIM XORCI_28 ( .CIN(\MUXCO_27|COUT_net ), .DIN(DX[28]), .SUM(
        SUM[28]) );
    CS_XORCI_PRIM XORCI_29 ( .CIN(\MUXCO_28|COUT_net ), .DIN(DX[29]), .SUM(
        SUM[29]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_30 ( .CIN(\MUXCO_29|COUT_net ), .DIN(DX[30]), .SUM(
        SUM[30]) );
    CS_XORCI_PRIM XORCI_31 ( .CIN(\MUXCO_30|COUT_net ), .DIN(DX[31]), .SUM(
        SUM[31]) );
    CS_XORCI_PRIM XORCI_32 ( .CIN(\MUXCO_31|COUT_net ), .DIN(DX[32]), .SUM(
        SUM[32]) );
    CS_XORCI_PRIM XORCI_33 ( .CIN(\MUXCO_32|COUT_net ), .DIN(DX[33]), .SUM(
        SUM[33]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
    CS_XORCI_PRIM XORCI_9 ( .CIN(\MUXCO_8|COUT_net ), .DIN(DX[9]), .SUM(SUM[9]) );
endmodule


module scaler_ipc_adder_7(CA, CI, CO, DX, SUM);
  input [6:0] CA;
  input CI;
  output CO;
  input [6:0] DX;
  output [6:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(CO), 
        .CSEL(DX[6]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
endmodule


module scaler_ipc_adder_8(CA, CI, CO, DX, SUM);
  input [7:0] CA;
  input CI;
  output CO;
  input [7:0] DX;
  output [7:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(CO), 
        .CSEL(DX[7]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
endmodule


module scaler_ipc_adder_9(CA, CI, CO, DX, SUM);
  input [8:0] CA;
  input CI;
  output CO;
  input [8:0] DX;
  output [8:0] SUM;

    wire \MUXCO_0|COUT_net ;
    wire \MUXCO_1|COUT_net ;
    wire \MUXCO_2|COUT_net ;
    wire \MUXCO_3|COUT_net ;
    wire \MUXCO_4|COUT_net ;
    wire \MUXCO_5|COUT_net ;
    wire \MUXCO_6|COUT_net ;
    wire \MUXCO_7|COUT_net ;

    CS_MUXCO_PRIM MUXCO_0 ( .AIN(CA[0]), .CIN(CI), .COUT(\MUXCO_0|COUT_net ), 
        .CSEL(DX[0]) );
    CS_MUXCO_PRIM MUXCO_1 ( .AIN(CA[1]), .CIN(\MUXCO_0|COUT_net ), .COUT(
        \MUXCO_1|COUT_net ), .CSEL(DX[1]) );
    CS_MUXCO_PRIM MUXCO_2 ( .AIN(CA[2]), .CIN(\MUXCO_1|COUT_net ), .COUT(
        \MUXCO_2|COUT_net ), .CSEL(DX[2]) );
    CS_MUXCO_PRIM MUXCO_3 ( .AIN(CA[3]), .CIN(\MUXCO_2|COUT_net ), .COUT(
        \MUXCO_3|COUT_net ), .CSEL(DX[3]) );
    CS_MUXCO_PRIM MUXCO_4 ( .AIN(CA[4]), .CIN(\MUXCO_3|COUT_net ), .COUT(
        \MUXCO_4|COUT_net ), .CSEL(DX[4]) );
    CS_MUXCO_PRIM MUXCO_5 ( .AIN(CA[5]), .CIN(\MUXCO_4|COUT_net ), .COUT(
        \MUXCO_5|COUT_net ), .CSEL(DX[5]) );
    CS_MUXCO_PRIM MUXCO_6 ( .AIN(CA[6]), .CIN(\MUXCO_5|COUT_net ), .COUT(
        \MUXCO_6|COUT_net ), .CSEL(DX[6]) );
    CS_MUXCO_PRIM MUXCO_7 ( .AIN(CA[7]), .CIN(\MUXCO_6|COUT_net ), .COUT(
        \MUXCO_7|COUT_net ), .CSEL(DX[7]) );
    CS_MUXCO_PRIM MUXCO_8 ( .AIN(CA[8]), .CIN(\MUXCO_7|COUT_net ), .COUT(CO), 
        .CSEL(DX[8]) );
    CS_XORCI_PRIM XORCI_0 ( .CIN(CI), .DIN(DX[0]), .SUM(SUM[0]) );
    CS_XORCI_PRIM XORCI_1 ( .CIN(\MUXCO_0|COUT_net ), .DIN(DX[1]), .SUM(SUM[1]) );
    CS_XORCI_PRIM XORCI_2 ( .CIN(\MUXCO_1|COUT_net ), .DIN(DX[2]), .SUM(SUM[2]) );
    CS_XORCI_PRIM XORCI_3 ( .CIN(\MUXCO_2|COUT_net ), .DIN(DX[3]), .SUM(SUM[3]) );
    CS_XORCI_PRIM XORCI_4 ( .CIN(\MUXCO_3|COUT_net ), .DIN(DX[4]), .SUM(SUM[4]) );
    CS_XORCI_PRIM XORCI_5 ( .CIN(\MUXCO_4|COUT_net ), .DIN(DX[5]), .SUM(SUM[5]) );
    CS_XORCI_PRIM XORCI_6 ( .CIN(\MUXCO_5|COUT_net ), .DIN(DX[6]), .SUM(SUM[6]) );
    CS_XORCI_PRIM XORCI_7 ( .CIN(\MUXCO_6|COUT_net ), .DIN(DX[7]), .SUM(SUM[7]) );
    CS_XORCI_PRIM XORCI_8 ( .CIN(\MUXCO_7|COUT_net ), .DIN(DX[8]), .SUM(SUM[8]) );
endmodule


module scaler ( HS, VS, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u138_mac, a_acc_en_cal1_u139_mac,
           a_acc_en_cal1_u140_mac, a_acc_en_cal1_u141_mac, a_acc_en_cal1_u142_mac,
           a_acc_en_cal1_u143_mac, a_acc_en_cal1_u144_mac, a_acc_en_cal1_u145_mac,
           a_acc_en_cal1_u146_mac, a_acc_en_cal1_u147_mac, a_acc_en_cal1_u148_mac,
           a_acc_en_cal1_u149_mac, a_acc_en_coefcal1_u63_mac, a_acc_en_coefcal1_u64_mac,
           a_acc_en_coefcal1_u64_mac_0_, \a_dinx[0]_cal1_u137_mac , \a_dinx[0]_cal1_u138_mac ,
           \a_dinx[0]_cal1_u139_mac , \a_dinx[0]_cal1_u140_mac , \a_dinx[0]_cal1_u141_mac ,
           \a_dinx[0]_cal1_u142_mac , \a_dinx[0]_cal1_u143_mac , \a_dinx[0]_cal1_u144_mac ,
           \a_dinx[0]_cal1_u145_mac , \a_dinx[0]_cal1_u146_mac , \a_dinx[0]_cal1_u147_mac ,
           \a_dinx[0]_cal1_u148_mac , \a_dinx[0]_cal1_u149_mac , \a_dinx[0]_coefcal1_u63_mac ,
           \a_dinx[0]_coefcal1_u64_mac , \a_dinx[0]_coefcal1_u64_mac_0_ ,
           \a_dinx[10]_cal1_u137_mac , \a_dinx[10]_cal1_u138_mac , \a_dinx[10]_cal1_u139_mac ,
           \a_dinx[10]_cal1_u140_mac , \a_dinx[10]_cal1_u141_mac , \a_dinx[10]_cal1_u142_mac ,
           \a_dinx[10]_cal1_u143_mac , \a_dinx[10]_cal1_u144_mac , \a_dinx[10]_cal1_u145_mac ,
           \a_dinx[10]_cal1_u146_mac , \a_dinx[10]_cal1_u147_mac , \a_dinx[10]_cal1_u148_mac ,
           \a_dinx[10]_cal1_u149_mac , \a_dinx[10]_coefcal1_u63_mac , \a_dinx[10]_coefcal1_u64_mac ,
           \a_dinx[10]_coefcal1_u64_mac_0_ , \a_dinx[11]_cal1_u137_mac , \a_dinx[11]_cal1_u138_mac ,
           \a_dinx[11]_cal1_u139_mac , \a_dinx[11]_cal1_u140_mac , \a_dinx[11]_cal1_u141_mac ,
           \a_dinx[11]_cal1_u142_mac , \a_dinx[11]_cal1_u143_mac , \a_dinx[11]_cal1_u144_mac ,
           \a_dinx[11]_cal1_u145_mac , \a_dinx[11]_cal1_u146_mac , \a_dinx[11]_cal1_u147_mac ,
           \a_dinx[11]_cal1_u148_mac , \a_dinx[11]_cal1_u149_mac , \a_dinx[11]_coefcal1_u63_mac ,
           \a_dinx[11]_coefcal1_u64_mac , \a_dinx[11]_coefcal1_u64_mac_0_ ,
           \a_dinx[12]_cal1_u137_mac , \a_dinx[12]_cal1_u138_mac , \a_dinx[12]_cal1_u139_mac ,
           \a_dinx[12]_cal1_u140_mac , \a_dinx[12]_cal1_u141_mac , \a_dinx[12]_cal1_u142_mac ,
           \a_dinx[12]_cal1_u143_mac , \a_dinx[12]_cal1_u144_mac , \a_dinx[12]_cal1_u145_mac ,
           \a_dinx[12]_cal1_u146_mac , \a_dinx[12]_cal1_u147_mac , \a_dinx[12]_cal1_u148_mac ,
           \a_dinx[12]_cal1_u149_mac , \a_dinx[12]_coefcal1_u63_mac , \a_dinx[12]_coefcal1_u64_mac ,
           \a_dinx[12]_coefcal1_u64_mac_0_ , \a_dinx[13]_cal1_u137_mac , \a_dinx[13]_cal1_u138_mac ,
           \a_dinx[13]_cal1_u139_mac , \a_dinx[13]_cal1_u140_mac , \a_dinx[13]_cal1_u141_mac ,
           \a_dinx[13]_cal1_u142_mac , \a_dinx[13]_cal1_u143_mac , \a_dinx[13]_cal1_u144_mac ,
           \a_dinx[13]_cal1_u145_mac , \a_dinx[13]_cal1_u146_mac , \a_dinx[13]_cal1_u147_mac ,
           \a_dinx[13]_cal1_u148_mac , \a_dinx[13]_cal1_u149_mac , \a_dinx[13]_coefcal1_u63_mac ,
           \a_dinx[13]_coefcal1_u64_mac , \a_dinx[13]_coefcal1_u64_mac_0_ ,
           \a_dinx[1]_cal1_u137_mac , \a_dinx[1]_cal1_u138_mac , \a_dinx[1]_cal1_u139_mac ,
           \a_dinx[1]_cal1_u140_mac , \a_dinx[1]_cal1_u141_mac , \a_dinx[1]_cal1_u142_mac ,
           \a_dinx[1]_cal1_u143_mac , \a_dinx[1]_cal1_u144_mac , \a_dinx[1]_cal1_u145_mac ,
           \a_dinx[1]_cal1_u146_mac , \a_dinx[1]_cal1_u147_mac , \a_dinx[1]_cal1_u148_mac ,
           \a_dinx[1]_cal1_u149_mac , \a_dinx[1]_coefcal1_u63_mac , \a_dinx[1]_coefcal1_u64_mac ,
           \a_dinx[1]_coefcal1_u64_mac_0_ , \a_dinx[2]_cal1_u137_mac , \a_dinx[2]_cal1_u138_mac ,
           \a_dinx[2]_cal1_u139_mac , \a_dinx[2]_cal1_u140_mac , \a_dinx[2]_cal1_u141_mac ,
           \a_dinx[2]_cal1_u142_mac , \a_dinx[2]_cal1_u143_mac , \a_dinx[2]_cal1_u144_mac ,
           \a_dinx[2]_cal1_u145_mac , \a_dinx[2]_cal1_u146_mac , \a_dinx[2]_cal1_u147_mac ,
           \a_dinx[2]_cal1_u148_mac , \a_dinx[2]_cal1_u149_mac , \a_dinx[2]_coefcal1_u63_mac ,
           \a_dinx[2]_coefcal1_u64_mac , \a_dinx[2]_coefcal1_u64_mac_0_ ,
           \a_dinx[3]_cal1_u137_mac , \a_dinx[3]_cal1_u138_mac , \a_dinx[3]_cal1_u139_mac ,
           \a_dinx[3]_cal1_u140_mac , \a_dinx[3]_cal1_u141_mac , \a_dinx[3]_cal1_u142_mac ,
           \a_dinx[3]_cal1_u143_mac , \a_dinx[3]_cal1_u144_mac , \a_dinx[3]_cal1_u145_mac ,
           \a_dinx[3]_cal1_u146_mac , \a_dinx[3]_cal1_u147_mac , \a_dinx[3]_cal1_u148_mac ,
           \a_dinx[3]_cal1_u149_mac , \a_dinx[3]_coefcal1_u63_mac , \a_dinx[3]_coefcal1_u64_mac ,
           \a_dinx[3]_coefcal1_u64_mac_0_ , \a_dinx[4]_cal1_u137_mac , \a_dinx[4]_cal1_u138_mac ,
           \a_dinx[4]_cal1_u139_mac , \a_dinx[4]_cal1_u140_mac , \a_dinx[4]_cal1_u141_mac ,
           \a_dinx[4]_cal1_u142_mac , \a_dinx[4]_cal1_u143_mac , \a_dinx[4]_cal1_u144_mac ,
           \a_dinx[4]_cal1_u145_mac , \a_dinx[4]_cal1_u146_mac , \a_dinx[4]_cal1_u147_mac ,
           \a_dinx[4]_cal1_u148_mac , \a_dinx[4]_cal1_u149_mac , \a_dinx[4]_coefcal1_u63_mac ,
           \a_dinx[4]_coefcal1_u64_mac , \a_dinx[4]_coefcal1_u64_mac_0_ ,
           \a_dinx[5]_cal1_u137_mac , \a_dinx[5]_cal1_u138_mac , \a_dinx[5]_cal1_u139_mac ,
           \a_dinx[5]_cal1_u140_mac , \a_dinx[5]_cal1_u141_mac , \a_dinx[5]_cal1_u142_mac ,
           \a_dinx[5]_cal1_u143_mac , \a_dinx[5]_cal1_u144_mac , \a_dinx[5]_cal1_u145_mac ,
           \a_dinx[5]_cal1_u146_mac , \a_dinx[5]_cal1_u147_mac , \a_dinx[5]_cal1_u148_mac ,
           \a_dinx[5]_cal1_u149_mac , \a_dinx[5]_coefcal1_u63_mac , \a_dinx[5]_coefcal1_u64_mac ,
           \a_dinx[5]_coefcal1_u64_mac_0_ , \a_dinx[6]_cal1_u137_mac , \a_dinx[6]_cal1_u138_mac ,
           \a_dinx[6]_cal1_u139_mac , \a_dinx[6]_cal1_u140_mac , \a_dinx[6]_cal1_u141_mac ,
           \a_dinx[6]_cal1_u142_mac , \a_dinx[6]_cal1_u143_mac , \a_dinx[6]_cal1_u144_mac ,
           \a_dinx[6]_cal1_u145_mac , \a_dinx[6]_cal1_u146_mac , \a_dinx[6]_cal1_u147_mac ,
           \a_dinx[6]_cal1_u148_mac , \a_dinx[6]_cal1_u149_mac , \a_dinx[6]_coefcal1_u63_mac ,
           \a_dinx[6]_coefcal1_u64_mac , \a_dinx[6]_coefcal1_u64_mac_0_ ,
           \a_dinx[7]_cal1_u137_mac , \a_dinx[7]_cal1_u138_mac , \a_dinx[7]_cal1_u139_mac ,
           \a_dinx[7]_cal1_u140_mac , \a_dinx[7]_cal1_u141_mac , \a_dinx[7]_cal1_u142_mac ,
           \a_dinx[7]_cal1_u143_mac , \a_dinx[7]_cal1_u144_mac , \a_dinx[7]_cal1_u145_mac ,
           \a_dinx[7]_cal1_u146_mac , \a_dinx[7]_cal1_u147_mac , \a_dinx[7]_cal1_u148_mac ,
           \a_dinx[7]_cal1_u149_mac , \a_dinx[7]_coefcal1_u63_mac , \a_dinx[7]_coefcal1_u64_mac ,
           \a_dinx[7]_coefcal1_u64_mac_0_ , \a_dinx[8]_cal1_u137_mac , \a_dinx[8]_cal1_u138_mac ,
           \a_dinx[8]_cal1_u139_mac , \a_dinx[8]_cal1_u140_mac , \a_dinx[8]_cal1_u141_mac ,
           \a_dinx[8]_cal1_u142_mac , \a_dinx[8]_cal1_u143_mac , \a_dinx[8]_cal1_u144_mac ,
           \a_dinx[8]_cal1_u145_mac , \a_dinx[8]_cal1_u146_mac , \a_dinx[8]_cal1_u147_mac ,
           \a_dinx[8]_cal1_u148_mac , \a_dinx[8]_cal1_u149_mac , \a_dinx[8]_coefcal1_u63_mac ,
           \a_dinx[8]_coefcal1_u64_mac , \a_dinx[8]_coefcal1_u64_mac_0_ ,
           \a_dinx[9]_cal1_u137_mac , \a_dinx[9]_cal1_u138_mac , \a_dinx[9]_cal1_u139_mac ,
           \a_dinx[9]_cal1_u140_mac , \a_dinx[9]_cal1_u141_mac , \a_dinx[9]_cal1_u142_mac ,
           \a_dinx[9]_cal1_u143_mac , \a_dinx[9]_cal1_u144_mac , \a_dinx[9]_cal1_u145_mac ,
           \a_dinx[9]_cal1_u146_mac , \a_dinx[9]_cal1_u147_mac , \a_dinx[9]_cal1_u148_mac ,
           \a_dinx[9]_cal1_u149_mac , \a_dinx[9]_coefcal1_u63_mac , \a_dinx[9]_coefcal1_u64_mac ,
           \a_dinx[9]_coefcal1_u64_mac_0_ , a_dinxy_cen_cal1_u137_mac, a_dinxy_cen_cal1_u138_mac,
           a_dinxy_cen_cal1_u139_mac, a_dinxy_cen_cal1_u140_mac, a_dinxy_cen_cal1_u141_mac,
           a_dinxy_cen_cal1_u142_mac, a_dinxy_cen_cal1_u143_mac, a_dinxy_cen_cal1_u144_mac,
           a_dinxy_cen_cal1_u145_mac, a_dinxy_cen_cal1_u146_mac, a_dinxy_cen_cal1_u147_mac,
           a_dinxy_cen_cal1_u148_mac, a_dinxy_cen_cal1_u149_mac, a_dinxy_cen_coefcal1_u63_mac,
           a_dinxy_cen_coefcal1_u64_mac, a_dinxy_cen_coefcal1_u64_mac_0_,
           \a_diny[0]_cal1_u137_mac , \a_diny[0]_cal1_u138_mac , \a_diny[0]_cal1_u139_mac ,
           \a_diny[0]_cal1_u140_mac , \a_diny[0]_cal1_u141_mac , \a_diny[0]_cal1_u142_mac ,
           \a_diny[0]_cal1_u143_mac , \a_diny[0]_cal1_u144_mac , \a_diny[0]_cal1_u145_mac ,
           \a_diny[0]_cal1_u146_mac , \a_diny[0]_cal1_u147_mac , \a_diny[0]_cal1_u148_mac ,
           \a_diny[0]_cal1_u149_mac , \a_diny[0]_coefcal1_u63_mac , \a_diny[0]_coefcal1_u64_mac ,
           \a_diny[0]_coefcal1_u64_mac_0_ , \a_diny[1]_cal1_u137_mac , \a_diny[1]_cal1_u138_mac ,
           \a_diny[1]_cal1_u139_mac , \a_diny[1]_cal1_u140_mac , \a_diny[1]_cal1_u141_mac ,
           \a_diny[1]_cal1_u142_mac , \a_diny[1]_cal1_u143_mac , \a_diny[1]_cal1_u144_mac ,
           \a_diny[1]_cal1_u145_mac , \a_diny[1]_cal1_u146_mac , \a_diny[1]_cal1_u147_mac ,
           \a_diny[1]_cal1_u148_mac , \a_diny[1]_cal1_u149_mac , \a_diny[1]_coefcal1_u63_mac ,
           \a_diny[1]_coefcal1_u64_mac , \a_diny[1]_coefcal1_u64_mac_0_ ,
           \a_diny[2]_cal1_u137_mac , \a_diny[2]_cal1_u138_mac , \a_diny[2]_cal1_u139_mac ,
           \a_diny[2]_cal1_u140_mac , \a_diny[2]_cal1_u141_mac , \a_diny[2]_cal1_u142_mac ,
           \a_diny[2]_cal1_u143_mac , \a_diny[2]_cal1_u144_mac , \a_diny[2]_cal1_u145_mac ,
           \a_diny[2]_cal1_u146_mac , \a_diny[2]_cal1_u147_mac , \a_diny[2]_cal1_u148_mac ,
           \a_diny[2]_cal1_u149_mac , \a_diny[2]_coefcal1_u63_mac , \a_diny[2]_coefcal1_u64_mac ,
           \a_diny[2]_coefcal1_u64_mac_0_ , \a_diny[3]_cal1_u137_mac , \a_diny[3]_cal1_u138_mac ,
           \a_diny[3]_cal1_u139_mac , \a_diny[3]_cal1_u140_mac , \a_diny[3]_cal1_u141_mac ,
           \a_diny[3]_cal1_u142_mac , \a_diny[3]_cal1_u143_mac , \a_diny[3]_cal1_u144_mac ,
           \a_diny[3]_cal1_u145_mac , \a_diny[3]_cal1_u146_mac , \a_diny[3]_cal1_u147_mac ,
           \a_diny[3]_cal1_u148_mac , \a_diny[3]_cal1_u149_mac , \a_diny[3]_coefcal1_u63_mac ,
           \a_diny[3]_coefcal1_u64_mac , \a_diny[3]_coefcal1_u64_mac_0_ ,
           \a_diny[4]_cal1_u137_mac , \a_diny[4]_cal1_u138_mac , \a_diny[4]_cal1_u139_mac ,
           \a_diny[4]_cal1_u140_mac , \a_diny[4]_cal1_u141_mac , \a_diny[4]_cal1_u142_mac ,
           \a_diny[4]_cal1_u143_mac , \a_diny[4]_cal1_u144_mac , \a_diny[4]_cal1_u145_mac ,
           \a_diny[4]_cal1_u146_mac , \a_diny[4]_cal1_u147_mac , \a_diny[4]_cal1_u148_mac ,
           \a_diny[4]_cal1_u149_mac , \a_diny[4]_coefcal1_u63_mac , \a_diny[4]_coefcal1_u64_mac ,
           \a_diny[4]_coefcal1_u64_mac_0_ , \a_diny[5]_cal1_u137_mac , \a_diny[5]_cal1_u138_mac ,
           \a_diny[5]_cal1_u139_mac , \a_diny[5]_cal1_u140_mac , \a_diny[5]_cal1_u141_mac ,
           \a_diny[5]_cal1_u142_mac , \a_diny[5]_cal1_u143_mac , \a_diny[5]_cal1_u144_mac ,
           \a_diny[5]_cal1_u145_mac , \a_diny[5]_cal1_u146_mac , \a_diny[5]_cal1_u147_mac ,
           \a_diny[5]_cal1_u148_mac , \a_diny[5]_cal1_u149_mac , \a_diny[5]_coefcal1_u63_mac ,
           \a_diny[5]_coefcal1_u64_mac , \a_diny[5]_coefcal1_u64_mac_0_ ,
           \a_diny[6]_cal1_u137_mac , \a_diny[6]_cal1_u138_mac , \a_diny[6]_cal1_u139_mac ,
           \a_diny[6]_cal1_u140_mac , \a_diny[6]_cal1_u141_mac , \a_diny[6]_cal1_u142_mac ,
           \a_diny[6]_cal1_u143_mac , \a_diny[6]_cal1_u144_mac , \a_diny[6]_cal1_u145_mac ,
           \a_diny[6]_cal1_u146_mac , \a_diny[6]_cal1_u147_mac , \a_diny[6]_cal1_u148_mac ,
           \a_diny[6]_cal1_u149_mac , \a_diny[6]_coefcal1_u63_mac , \a_diny[6]_coefcal1_u64_mac ,
           \a_diny[6]_coefcal1_u64_mac_0_ , \a_diny[7]_cal1_u137_mac , \a_diny[7]_cal1_u138_mac ,
           \a_diny[7]_cal1_u139_mac , \a_diny[7]_cal1_u140_mac , \a_diny[7]_cal1_u141_mac ,
           \a_diny[7]_cal1_u142_mac , \a_diny[7]_cal1_u143_mac , \a_diny[7]_cal1_u144_mac ,
           \a_diny[7]_cal1_u145_mac , \a_diny[7]_cal1_u146_mac , \a_diny[7]_cal1_u147_mac ,
           \a_diny[7]_cal1_u148_mac , \a_diny[7]_cal1_u149_mac , \a_diny[7]_coefcal1_u63_mac ,
           \a_diny[7]_coefcal1_u64_mac , \a_diny[7]_coefcal1_u64_mac_0_ ,
           \a_diny[8]_cal1_u137_mac , \a_diny[8]_cal1_u138_mac , \a_diny[8]_cal1_u139_mac ,
           \a_diny[8]_cal1_u140_mac , \a_diny[8]_cal1_u141_mac , \a_diny[8]_cal1_u142_mac ,
           \a_diny[8]_cal1_u143_mac , \a_diny[8]_cal1_u144_mac , \a_diny[8]_cal1_u145_mac ,
           \a_diny[8]_cal1_u146_mac , \a_diny[8]_cal1_u147_mac , \a_diny[8]_cal1_u148_mac ,
           \a_diny[8]_cal1_u149_mac , \a_diny[8]_coefcal1_u63_mac , \a_diny[8]_coefcal1_u64_mac ,
           \a_diny[8]_coefcal1_u64_mac_0_ , \a_diny[9]_cal1_u137_mac , \a_diny[9]_cal1_u138_mac ,
           \a_diny[9]_cal1_u139_mac , \a_diny[9]_cal1_u140_mac , \a_diny[9]_cal1_u141_mac ,
           \a_diny[9]_cal1_u142_mac , \a_diny[9]_cal1_u143_mac , \a_diny[9]_cal1_u144_mac ,
           \a_diny[9]_cal1_u145_mac , \a_diny[9]_cal1_u146_mac , \a_diny[9]_cal1_u147_mac ,
           \a_diny[9]_cal1_u148_mac , \a_diny[9]_cal1_u149_mac , \a_diny[9]_coefcal1_u63_mac ,
           \a_diny[9]_coefcal1_u64_mac , \a_diny[9]_coefcal1_u64_mac_0_ ,
           a_dinz_cen_cal1_u137_mac, a_dinz_cen_cal1_u138_mac, a_dinz_cen_cal1_u139_mac,
           a_dinz_cen_cal1_u140_mac, a_dinz_cen_cal1_u141_mac, a_dinz_cen_cal1_u142_mac,
           a_dinz_cen_cal1_u143_mac, a_dinz_cen_cal1_u144_mac, a_dinz_cen_cal1_u145_mac,
           a_dinz_cen_cal1_u146_mac, a_dinz_cen_cal1_u147_mac, a_dinz_cen_cal1_u148_mac,
           a_dinz_cen_cal1_u149_mac, a_dinz_cen_coefcal1_u63_mac, a_dinz_cen_coefcal1_u64_mac,
           a_dinz_cen_coefcal1_u64_mac_0_, a_dinz_en_cal1_u137_mac, a_dinz_en_cal1_u138_mac,
           a_dinz_en_cal1_u139_mac, a_dinz_en_cal1_u140_mac, a_dinz_en_cal1_u141_mac,
           a_dinz_en_cal1_u142_mac, a_dinz_en_cal1_u143_mac, a_dinz_en_cal1_u144_mac,
           a_dinz_en_cal1_u145_mac, a_dinz_en_cal1_u146_mac, a_dinz_en_cal1_u147_mac,
           a_dinz_en_cal1_u148_mac, a_dinz_en_cal1_u149_mac, a_dinz_en_coefcal1_u63_mac,
           a_dinz_en_coefcal1_u64_mac, a_dinz_en_coefcal1_u64_mac_0_, a_in_sr_cal1_u137_mac,
           a_in_sr_cal1_u138_mac, a_in_sr_cal1_u139_mac, a_in_sr_cal1_u140_mac,
           a_in_sr_cal1_u141_mac, a_in_sr_cal1_u142_mac, a_in_sr_cal1_u143_mac,
           a_in_sr_cal1_u144_mac, a_in_sr_cal1_u145_mac, a_in_sr_cal1_u146_mac,
           a_in_sr_cal1_u147_mac, a_in_sr_cal1_u148_mac, a_in_sr_cal1_u149_mac,
           a_in_sr_coefcal1_u63_mac, a_in_sr_coefcal1_u64_mac, a_in_sr_coefcal1_u64_mac_0_,
           \a_mac_out[0]_coefcal1_u63_mac , \a_mac_out[0]_coefcal1_u64_mac ,
           \a_mac_out[0]_coefcal1_u64_mac_0_ , \a_mac_out[10]_cal1_u137_mac ,
           \a_mac_out[10]_cal1_u138_mac , \a_mac_out[10]_cal1_u139_mac , \a_mac_out[10]_cal1_u140_mac ,
           \a_mac_out[10]_cal1_u141_mac , \a_mac_out[10]_cal1_u142_mac , \a_mac_out[10]_cal1_u143_mac ,
           \a_mac_out[10]_cal1_u144_mac , \a_mac_out[10]_cal1_u145_mac , \a_mac_out[10]_cal1_u146_mac ,
           \a_mac_out[10]_cal1_u147_mac , \a_mac_out[10]_cal1_u148_mac , \a_mac_out[10]_cal1_u149_mac ,
           \a_mac_out[10]_coefcal1_u63_mac , \a_mac_out[10]_coefcal1_u64_mac ,
           \a_mac_out[10]_coefcal1_u64_mac_0_ , \a_mac_out[11]_cal1_u137_mac ,
           \a_mac_out[11]_cal1_u138_mac , \a_mac_out[11]_cal1_u139_mac , \a_mac_out[11]_cal1_u140_mac ,
           \a_mac_out[11]_cal1_u141_mac , \a_mac_out[11]_cal1_u142_mac , \a_mac_out[11]_cal1_u143_mac ,
           \a_mac_out[11]_cal1_u144_mac , \a_mac_out[11]_cal1_u145_mac , \a_mac_out[11]_cal1_u146_mac ,
           \a_mac_out[11]_cal1_u147_mac , \a_mac_out[11]_cal1_u148_mac , \a_mac_out[11]_cal1_u149_mac ,
           \a_mac_out[11]_coefcal1_u63_mac , \a_mac_out[11]_coefcal1_u64_mac ,
           \a_mac_out[11]_coefcal1_u64_mac_0_ , \a_mac_out[12]_cal1_u138_mac ,
           \a_mac_out[12]_cal1_u139_mac , \a_mac_out[12]_cal1_u140_mac , \a_mac_out[12]_cal1_u141_mac ,
           \a_mac_out[12]_cal1_u142_mac , \a_mac_out[12]_cal1_u143_mac , \a_mac_out[12]_cal1_u144_mac ,
           \a_mac_out[12]_cal1_u145_mac , \a_mac_out[12]_cal1_u146_mac , \a_mac_out[12]_cal1_u147_mac ,
           \a_mac_out[12]_cal1_u148_mac , \a_mac_out[12]_cal1_u149_mac , \a_mac_out[12]_coefcal1_u63_mac ,
           \a_mac_out[12]_coefcal1_u64_mac , \a_mac_out[12]_coefcal1_u64_mac_0_ ,
           \a_mac_out[13]_cal1_u138_mac , \a_mac_out[13]_cal1_u139_mac , \a_mac_out[13]_cal1_u140_mac ,
           \a_mac_out[13]_cal1_u141_mac , \a_mac_out[13]_cal1_u142_mac , \a_mac_out[13]_cal1_u143_mac ,
           \a_mac_out[13]_cal1_u144_mac , \a_mac_out[13]_cal1_u145_mac , \a_mac_out[13]_cal1_u146_mac ,
           \a_mac_out[13]_cal1_u147_mac , \a_mac_out[13]_cal1_u148_mac , \a_mac_out[13]_cal1_u149_mac ,
           \a_mac_out[13]_coefcal1_u63_mac , \a_mac_out[13]_coefcal1_u64_mac ,
           \a_mac_out[14]_coefcal1_u63_mac , \a_mac_out[14]_coefcal1_u64_mac ,
           \a_mac_out[15]_coefcal1_u63_mac , \a_mac_out[15]_coefcal1_u64_mac ,
           \a_mac_out[16]_coefcal1_u63_mac , \a_mac_out[16]_coefcal1_u64_mac ,
           \a_mac_out[17]_coefcal1_u63_mac , \a_mac_out[17]_coefcal1_u64_mac ,
           \a_mac_out[18]_coefcal1_u63_mac , \a_mac_out[18]_coefcal1_u64_mac ,
           \a_mac_out[19]_coefcal1_u63_mac , \a_mac_out[19]_coefcal1_u64_mac ,
           \a_mac_out[1]_coefcal1_u63_mac , \a_mac_out[1]_coefcal1_u64_mac ,
           \a_mac_out[1]_coefcal1_u64_mac_0_ , \a_mac_out[20]_coefcal1_u64_mac ,
           \a_mac_out[21]_coefcal1_u64_mac , \a_mac_out[22]_coefcal1_u64_mac ,
           \a_mac_out[23]_coefcal1_u64_mac , \a_mac_out[2]_coefcal1_u63_mac ,
           \a_mac_out[2]_coefcal1_u64_mac , \a_mac_out[2]_coefcal1_u64_mac_0_ ,
           \a_mac_out[3]_coefcal1_u63_mac , \a_mac_out[3]_coefcal1_u64_mac ,
           \a_mac_out[3]_coefcal1_u64_mac_0_ , \a_mac_out[4]_coefcal1_u63_mac ,
           \a_mac_out[4]_coefcal1_u64_mac , \a_mac_out[4]_coefcal1_u64_mac_0_ ,
           \a_mac_out[5]_coefcal1_u63_mac , \a_mac_out[5]_coefcal1_u64_mac ,
           \a_mac_out[5]_coefcal1_u64_mac_0_ , \a_mac_out[6]_cal1_u137_mac ,
           \a_mac_out[6]_cal1_u138_mac , \a_mac_out[6]_cal1_u139_mac , \a_mac_out[6]_cal1_u140_mac ,
           \a_mac_out[6]_cal1_u141_mac , \a_mac_out[6]_cal1_u142_mac , \a_mac_out[6]_cal1_u143_mac ,
           \a_mac_out[6]_cal1_u144_mac , \a_mac_out[6]_cal1_u145_mac , \a_mac_out[6]_cal1_u146_mac ,
           \a_mac_out[6]_cal1_u147_mac , \a_mac_out[6]_cal1_u148_mac , \a_mac_out[6]_cal1_u149_mac ,
           \a_mac_out[6]_coefcal1_u63_mac , \a_mac_out[6]_coefcal1_u64_mac ,
           \a_mac_out[6]_coefcal1_u64_mac_0_ , \a_mac_out[7]_cal1_u137_mac ,
           \a_mac_out[7]_cal1_u138_mac , \a_mac_out[7]_cal1_u139_mac , \a_mac_out[7]_cal1_u140_mac ,
           \a_mac_out[7]_cal1_u141_mac , \a_mac_out[7]_cal1_u142_mac , \a_mac_out[7]_cal1_u143_mac ,
           \a_mac_out[7]_cal1_u144_mac , \a_mac_out[7]_cal1_u145_mac , \a_mac_out[7]_cal1_u146_mac ,
           \a_mac_out[7]_cal1_u147_mac , \a_mac_out[7]_cal1_u148_mac , \a_mac_out[7]_cal1_u149_mac ,
           \a_mac_out[7]_coefcal1_u63_mac , \a_mac_out[7]_coefcal1_u64_mac ,
           \a_mac_out[7]_coefcal1_u64_mac_0_ , \a_mac_out[8]_cal1_u137_mac ,
           \a_mac_out[8]_cal1_u138_mac , \a_mac_out[8]_cal1_u139_mac , \a_mac_out[8]_cal1_u140_mac ,
           \a_mac_out[8]_cal1_u141_mac , \a_mac_out[8]_cal1_u142_mac , \a_mac_out[8]_cal1_u143_mac ,
           \a_mac_out[8]_cal1_u144_mac , \a_mac_out[8]_cal1_u145_mac , \a_mac_out[8]_cal1_u146_mac ,
           \a_mac_out[8]_cal1_u147_mac , \a_mac_out[8]_cal1_u148_mac , \a_mac_out[8]_cal1_u149_mac ,
           \a_mac_out[8]_coefcal1_u63_mac , \a_mac_out[8]_coefcal1_u64_mac ,
           \a_mac_out[8]_coefcal1_u64_mac_0_ , \a_mac_out[9]_cal1_u137_mac ,
           \a_mac_out[9]_cal1_u138_mac , \a_mac_out[9]_cal1_u139_mac , \a_mac_out[9]_cal1_u140_mac ,
           \a_mac_out[9]_cal1_u141_mac , \a_mac_out[9]_cal1_u142_mac , \a_mac_out[9]_cal1_u143_mac ,
           \a_mac_out[9]_cal1_u144_mac , \a_mac_out[9]_cal1_u145_mac , \a_mac_out[9]_cal1_u146_mac ,
           \a_mac_out[9]_cal1_u147_mac , \a_mac_out[9]_cal1_u148_mac , \a_mac_out[9]_cal1_u149_mac ,
           \a_mac_out[9]_coefcal1_u63_mac , \a_mac_out[9]_coefcal1_u64_mac ,
           \a_mac_out[9]_coefcal1_u64_mac_0_ , a_mac_out_cen_cal1_u137_mac,
           a_mac_out_cen_cal1_u138_mac, a_mac_out_cen_cal1_u139_mac, a_mac_out_cen_cal1_u140_mac,
           a_mac_out_cen_cal1_u141_mac, a_mac_out_cen_cal1_u142_mac, a_mac_out_cen_cal1_u143_mac,
           a_mac_out_cen_cal1_u144_mac, a_mac_out_cen_cal1_u145_mac, a_mac_out_cen_cal1_u146_mac,
           a_mac_out_cen_cal1_u147_mac, a_mac_out_cen_cal1_u148_mac, a_mac_out_cen_cal1_u149_mac,
           a_mac_out_cen_coefcal1_u63_mac, a_mac_out_cen_coefcal1_u64_mac,
           a_mac_out_cen_coefcal1_u64_mac_0_, a_out_sr_cal1_u137_mac, a_out_sr_cal1_u138_mac,
           a_out_sr_cal1_u139_mac, a_out_sr_cal1_u140_mac, a_out_sr_cal1_u141_mac,
           a_out_sr_cal1_u142_mac, a_out_sr_cal1_u143_mac, a_out_sr_cal1_u144_mac,
           a_out_sr_cal1_u145_mac, a_out_sr_cal1_u146_mac, a_out_sr_cal1_u147_mac,
           a_out_sr_cal1_u148_mac, a_out_sr_cal1_u149_mac, a_out_sr_coefcal1_u63_mac,
           a_out_sr_coefcal1_u64_mac, a_out_sr_coefcal1_u64_mac_0_, a_sload_cal1_u137_mac,
           a_sload_cal1_u138_mac, a_sload_cal1_u139_mac, a_sload_cal1_u140_mac,
           a_sload_cal1_u141_mac, a_sload_cal1_u142_mac, a_sload_cal1_u143_mac,
           a_sload_cal1_u144_mac, a_sload_cal1_u145_mac, a_sload_cal1_u146_mac,
           a_sload_cal1_u147_mac, a_sload_cal1_u148_mac, a_sload_cal1_u149_mac,
           a_sload_coefcal1_u63_mac, a_sload_coefcal1_u64_mac, a_sload_coefcal1_u64_mac_0_,
           b_acc_en_coefcal1_u64_mac, b_acc_en_coefcal1_u64_mac_0_, \b_dinx[0]_coefcal1_u64_mac ,
           \b_dinx[0]_coefcal1_u64_mac_0_ , \b_dinx[10]_coefcal1_u64_mac ,
           \b_dinx[10]_coefcal1_u64_mac_0_ , \b_dinx[11]_coefcal1_u64_mac ,
           \b_dinx[11]_coefcal1_u64_mac_0_ , \b_dinx[12]_coefcal1_u64_mac ,
           \b_dinx[12]_coefcal1_u64_mac_0_ , \b_dinx[13]_coefcal1_u64_mac ,
           \b_dinx[13]_coefcal1_u64_mac_0_ , \b_dinx[1]_coefcal1_u64_mac ,
           \b_dinx[1]_coefcal1_u64_mac_0_ , \b_dinx[2]_coefcal1_u64_mac ,
           \b_dinx[2]_coefcal1_u64_mac_0_ , \b_dinx[3]_coefcal1_u64_mac ,
           \b_dinx[3]_coefcal1_u64_mac_0_ , \b_dinx[4]_coefcal1_u64_mac ,
           \b_dinx[4]_coefcal1_u64_mac_0_ , \b_dinx[5]_coefcal1_u64_mac ,
           \b_dinx[5]_coefcal1_u64_mac_0_ , \b_dinx[6]_coefcal1_u64_mac ,
           \b_dinx[6]_coefcal1_u64_mac_0_ , \b_dinx[7]_coefcal1_u64_mac ,
           \b_dinx[7]_coefcal1_u64_mac_0_ , \b_dinx[8]_coefcal1_u64_mac ,
           \b_dinx[8]_coefcal1_u64_mac_0_ , \b_dinx[9]_coefcal1_u64_mac ,
           \b_dinx[9]_coefcal1_u64_mac_0_ , b_dinxy_cen_coefcal1_u64_mac,
           b_dinxy_cen_coefcal1_u64_mac_0_, \b_diny[0]_coefcal1_u64_mac ,
           \b_diny[0]_coefcal1_u64_mac_0_ , \b_diny[1]_coefcal1_u64_mac ,
           \b_diny[1]_coefcal1_u64_mac_0_ , \b_diny[2]_coefcal1_u64_mac ,
           \b_diny[2]_coefcal1_u64_mac_0_ , \b_diny[3]_coefcal1_u64_mac ,
           \b_diny[3]_coefcal1_u64_mac_0_ , \b_diny[4]_coefcal1_u64_mac ,
           \b_diny[4]_coefcal1_u64_mac_0_ , \b_diny[5]_coefcal1_u64_mac ,
           \b_diny[5]_coefcal1_u64_mac_0_ , \b_diny[6]_coefcal1_u64_mac ,
           \b_diny[6]_coefcal1_u64_mac_0_ , \b_diny[7]_coefcal1_u64_mac ,
           \b_diny[7]_coefcal1_u64_mac_0_ , \b_diny[8]_coefcal1_u64_mac ,
           \b_diny[8]_coefcal1_u64_mac_0_ , \b_diny[9]_coefcal1_u64_mac ,
           \b_diny[9]_coefcal1_u64_mac_0_ , b_dinz_cen_coefcal1_u64_mac, b_dinz_cen_coefcal1_u64_mac_0_,
           b_dinz_en_coefcal1_u64_mac, b_dinz_en_coefcal1_u64_mac_0_, b_in_sr_coefcal1_u64_mac,
           b_in_sr_coefcal1_u64_mac_0_, \b_mac_out[0]_coefcal1_u64_mac , \b_mac_out[1]_coefcal1_u64_mac ,
           \b_mac_out[2]_coefcal1_u64_mac , \b_mac_out[3]_coefcal1_u64_mac ,
           \b_mac_out[4]_coefcal1_u64_mac , b_mac_out_cen_coefcal1_u64_mac,
           b_mac_out_cen_coefcal1_u64_mac_0_, b_out_sr_coefcal1_u64_mac, b_out_sr_coefcal1_u64_mac_0_,
           b_sload_coefcal1_u64_mac, b_sload_coefcal1_u64_mac_0_, \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_1 , c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_0A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_0B_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_0B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_1A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1B_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_1B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2A_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_2A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2B_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_2B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3A_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_3A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3B_u_emb18k_0,
           c1r1_clka_fifo1_ram_inst_3B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_1, \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_q[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r1_q[9]_fifo1_ram_inst_3B_u_emb18k_1 , c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_1, c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_0,
           c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_1, c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_1, c1r2_clka_fifo1_ram_inst_0A_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_0A_u_emb18k_1, c1r2_clka_fifo1_ram_inst_0B_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_0B_u_emb18k_1, c1r2_clka_fifo1_ram_inst_1A_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_1A_u_emb18k_1, c1r2_clka_fifo1_ram_inst_1B_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_1B_u_emb18k_1, c1r2_clka_fifo1_ram_inst_2A_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_2A_u_emb18k_1, c1r2_clka_fifo1_ram_inst_2B_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_2B_u_emb18k_1, c1r2_clka_fifo1_ram_inst_3A_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_3A_u_emb18k_1, c1r2_clka_fifo1_ram_inst_3B_u_emb18k_0,
           c1r2_clka_fifo1_ram_inst_3B_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_1, c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_1, \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r2_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r2_q[9]_fifo1_ram_inst_3B_u_emb18k_0 , c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_1, c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_0,
           c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_1, c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_1, c1r3_clka_fifo1_ram_inst_0A_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_0A_u_emb18k_1, c1r3_clka_fifo1_ram_inst_0B_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_0B_u_emb18k_1, c1r3_clka_fifo1_ram_inst_1A_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_1A_u_emb18k_1, c1r3_clka_fifo1_ram_inst_1B_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_1B_u_emb18k_1, c1r3_clka_fifo1_ram_inst_2A_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_2A_u_emb18k_1, c1r3_clka_fifo1_ram_inst_2B_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_2B_u_emb18k_1, c1r3_clka_fifo1_ram_inst_3A_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_3A_u_emb18k_1, c1r3_clka_fifo1_ram_inst_3B_u_emb18k_0,
           c1r3_clka_fifo1_ram_inst_3B_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_1, c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_1, \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r3_q[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r3_q[9]_fifo1_ram_inst_3B_u_emb18k_1 , c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_1, c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_0,
           c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_1, c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_1, c1r4_clka_fifo1_ram_inst_0A_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_0A_u_emb18k_1, c1r4_clka_fifo1_ram_inst_0B_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_0B_u_emb18k_1, c1r4_clka_fifo1_ram_inst_1A_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_1A_u_emb18k_1, c1r4_clka_fifo1_ram_inst_1B_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_1B_u_emb18k_1, c1r4_clka_fifo1_ram_inst_2A_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_2A_u_emb18k_1, c1r4_clka_fifo1_ram_inst_2B_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_2B_u_emb18k_1, c1r4_clka_fifo1_ram_inst_3A_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_3A_u_emb18k_1, c1r4_clka_fifo1_ram_inst_3B_u_emb18k_0,
           c1r4_clka_fifo1_ram_inst_3B_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_1, c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_1, \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
           \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r4_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
           \c1r4_q[9]_fifo1_ram_inst_3B_u_emb18k_0 , c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_1, c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_0,
           c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_1, c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_0,
           c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_1, cea_fifo1_ram_inst_0A_u_emb18k_0,
           cea_fifo1_ram_inst_0A_u_emb18k_1, cea_fifo1_ram_inst_0B_u_emb18k_0,
           cea_fifo1_ram_inst_0B_u_emb18k_1, cea_fifo1_ram_inst_1A_u_emb18k_0,
           cea_fifo1_ram_inst_1A_u_emb18k_1, cea_fifo1_ram_inst_1B_u_emb18k_0,
           cea_fifo1_ram_inst_1B_u_emb18k_1, cea_fifo1_ram_inst_2A_u_emb18k_0,
           cea_fifo1_ram_inst_2A_u_emb18k_1, cea_fifo1_ram_inst_2B_u_emb18k_0,
           cea_fifo1_ram_inst_2B_u_emb18k_1, cea_fifo1_ram_inst_3A_u_emb18k_0,
           cea_fifo1_ram_inst_3A_u_emb18k_1, cea_fifo1_ram_inst_3B_u_emb18k_0,
           cea_fifo1_ram_inst_3B_u_emb18k_1, ceb_fifo1_ram_inst_0A_u_emb18k_0,
           ceb_fifo1_ram_inst_0A_u_emb18k_1, ceb_fifo1_ram_inst_0B_u_emb18k_0,
           ceb_fifo1_ram_inst_0B_u_emb18k_1, ceb_fifo1_ram_inst_1A_u_emb18k_0,
           ceb_fifo1_ram_inst_1A_u_emb18k_1, ceb_fifo1_ram_inst_1B_u_emb18k_0,
           ceb_fifo1_ram_inst_1B_u_emb18k_1, ceb_fifo1_ram_inst_2A_u_emb18k_0,
           ceb_fifo1_ram_inst_2A_u_emb18k_1, ceb_fifo1_ram_inst_2B_u_emb18k_0,
           ceb_fifo1_ram_inst_2B_u_emb18k_1, ceb_fifo1_ram_inst_3A_u_emb18k_0,
           ceb_fifo1_ram_inst_3A_u_emb18k_1, ceb_fifo1_ram_inst_3B_u_emb18k_0,
           ceb_fifo1_ram_inst_3B_u_emb18k_1, clka, clkb, dIn, dInEn, dOut,
           dOutEn, en, \haa[0]_fifo1_ram_inst_0A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_0B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_1B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_2A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_2B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_3A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
           \haa[0]_fifo1_ram_inst_3B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_0A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_0B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_1A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_1B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_2A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_2B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_3A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
           \haa[1]_fifo1_ram_inst_3B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_0A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_0B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_1A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_1B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_2A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_2B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_3A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
           \hab[0]_fifo1_ram_inst_3B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_0A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_0B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_1A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_1B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_2A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_2B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_3A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
           \hab[1]_fifo1_ram_inst_3B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
           iHsyn, iVsyn, inXRes, inYRes, outXRes, outYRes, rst, u5018_OUT,
           u5502_I1, u5502_I1_5_, u5502_IN, u5859_I1, u8205_O, u8205_O_1_,
           u8205_O_2_, u8218_Y, u8224_O, u8224_O_4_, u8230_O, u8231_O, u8245_D0,
           u8245_I0, u8245_I0_0_, u8245_I0_3_, u8245_IN, wea_fifo1_ram_inst_0A_u_emb18k_0,
           wea_fifo1_ram_inst_0A_u_emb18k_1, wea_fifo1_ram_inst_0B_u_emb18k_0,
           wea_fifo1_ram_inst_0B_u_emb18k_1, wea_fifo1_ram_inst_1A_u_emb18k_0,
           wea_fifo1_ram_inst_1A_u_emb18k_1, wea_fifo1_ram_inst_1B_u_emb18k_0,
           wea_fifo1_ram_inst_1B_u_emb18k_1, wea_fifo1_ram_inst_2A_u_emb18k_0,
           wea_fifo1_ram_inst_2A_u_emb18k_1, wea_fifo1_ram_inst_2B_u_emb18k_0,
           wea_fifo1_ram_inst_2B_u_emb18k_1, wea_fifo1_ram_inst_3A_u_emb18k_0,
           wea_fifo1_ram_inst_3A_u_emb18k_1, wea_fifo1_ram_inst_3B_u_emb18k_0,
           wea_fifo1_ram_inst_3B_u_emb18k_1, web_fifo1_ram_inst_0A_u_emb18k_0,
           web_fifo1_ram_inst_0A_u_emb18k_1, web_fifo1_ram_inst_0B_u_emb18k_0,
           web_fifo1_ram_inst_0B_u_emb18k_1, web_fifo1_ram_inst_1A_u_emb18k_0,
           web_fifo1_ram_inst_1A_u_emb18k_1, web_fifo1_ram_inst_1B_u_emb18k_0,
           web_fifo1_ram_inst_1B_u_emb18k_1, web_fifo1_ram_inst_2A_u_emb18k_0,
           web_fifo1_ram_inst_2A_u_emb18k_1, web_fifo1_ram_inst_2B_u_emb18k_0,
           web_fifo1_ram_inst_2B_u_emb18k_1, web_fifo1_ram_inst_3A_u_emb18k_0,
           web_fifo1_ram_inst_3A_u_emb18k_1, web_fifo1_ram_inst_3B_u_emb18k_0,
           web_fifo1_ram_inst_3B_u_emb18k_1, xBgn, xEnd, yBgn, yEnd );

    output HS, VS, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u138_mac, a_acc_en_cal1_u139_mac,
       a_acc_en_cal1_u140_mac, a_acc_en_cal1_u141_mac, a_acc_en_cal1_u142_mac,
       a_acc_en_cal1_u143_mac, a_acc_en_cal1_u144_mac, a_acc_en_cal1_u145_mac,
       a_acc_en_cal1_u146_mac, a_acc_en_cal1_u147_mac, a_acc_en_cal1_u148_mac,
       a_acc_en_cal1_u149_mac, a_acc_en_coefcal1_u63_mac, a_acc_en_coefcal1_u64_mac,
       a_acc_en_coefcal1_u64_mac_0_, \a_dinx[0]_cal1_u137_mac , \a_dinx[0]_cal1_u138_mac ,
       \a_dinx[0]_cal1_u139_mac , \a_dinx[0]_cal1_u140_mac , \a_dinx[0]_cal1_u141_mac ,
       \a_dinx[0]_cal1_u142_mac , \a_dinx[0]_cal1_u143_mac , \a_dinx[0]_cal1_u144_mac ,
       \a_dinx[0]_cal1_u145_mac , \a_dinx[0]_cal1_u146_mac , \a_dinx[0]_cal1_u147_mac ,
       \a_dinx[0]_cal1_u148_mac , \a_dinx[0]_cal1_u149_mac , \a_dinx[0]_coefcal1_u63_mac ,
       \a_dinx[0]_coefcal1_u64_mac , \a_dinx[0]_coefcal1_u64_mac_0_ , \a_dinx[10]_cal1_u137_mac ,
       \a_dinx[10]_cal1_u138_mac , \a_dinx[10]_cal1_u139_mac , \a_dinx[10]_cal1_u140_mac ,
       \a_dinx[10]_cal1_u141_mac , \a_dinx[10]_cal1_u142_mac , \a_dinx[10]_cal1_u143_mac ,
       \a_dinx[10]_cal1_u144_mac , \a_dinx[10]_cal1_u145_mac , \a_dinx[10]_cal1_u146_mac ,
       \a_dinx[10]_cal1_u147_mac , \a_dinx[10]_cal1_u148_mac , \a_dinx[10]_cal1_u149_mac ,
       \a_dinx[10]_coefcal1_u63_mac , \a_dinx[10]_coefcal1_u64_mac , \a_dinx[10]_coefcal1_u64_mac_0_ ,
       \a_dinx[11]_cal1_u137_mac , \a_dinx[11]_cal1_u138_mac , \a_dinx[11]_cal1_u139_mac ,
       \a_dinx[11]_cal1_u140_mac , \a_dinx[11]_cal1_u141_mac , \a_dinx[11]_cal1_u142_mac ,
       \a_dinx[11]_cal1_u143_mac , \a_dinx[11]_cal1_u144_mac , \a_dinx[11]_cal1_u145_mac ,
       \a_dinx[11]_cal1_u146_mac , \a_dinx[11]_cal1_u147_mac , \a_dinx[11]_cal1_u148_mac ,
       \a_dinx[11]_cal1_u149_mac , \a_dinx[11]_coefcal1_u63_mac , \a_dinx[11]_coefcal1_u64_mac ,
       \a_dinx[11]_coefcal1_u64_mac_0_ , \a_dinx[12]_cal1_u137_mac , \a_dinx[12]_cal1_u138_mac ,
       \a_dinx[12]_cal1_u139_mac , \a_dinx[12]_cal1_u140_mac , \a_dinx[12]_cal1_u141_mac ,
       \a_dinx[12]_cal1_u142_mac , \a_dinx[12]_cal1_u143_mac , \a_dinx[12]_cal1_u144_mac ,
       \a_dinx[12]_cal1_u145_mac , \a_dinx[12]_cal1_u146_mac , \a_dinx[12]_cal1_u147_mac ,
       \a_dinx[12]_cal1_u148_mac , \a_dinx[12]_cal1_u149_mac , \a_dinx[12]_coefcal1_u63_mac ,
       \a_dinx[12]_coefcal1_u64_mac , \a_dinx[12]_coefcal1_u64_mac_0_ , \a_dinx[13]_cal1_u137_mac ,
       \a_dinx[13]_cal1_u138_mac , \a_dinx[13]_cal1_u139_mac , \a_dinx[13]_cal1_u140_mac ,
       \a_dinx[13]_cal1_u141_mac , \a_dinx[13]_cal1_u142_mac , \a_dinx[13]_cal1_u143_mac ,
       \a_dinx[13]_cal1_u144_mac , \a_dinx[13]_cal1_u145_mac , \a_dinx[13]_cal1_u146_mac ,
       \a_dinx[13]_cal1_u147_mac , \a_dinx[13]_cal1_u148_mac , \a_dinx[13]_cal1_u149_mac ,
       \a_dinx[13]_coefcal1_u63_mac , \a_dinx[13]_coefcal1_u64_mac , \a_dinx[13]_coefcal1_u64_mac_0_ ,
       \a_dinx[1]_cal1_u137_mac , \a_dinx[1]_cal1_u138_mac , \a_dinx[1]_cal1_u139_mac ,
       \a_dinx[1]_cal1_u140_mac , \a_dinx[1]_cal1_u141_mac , \a_dinx[1]_cal1_u142_mac ,
       \a_dinx[1]_cal1_u143_mac , \a_dinx[1]_cal1_u144_mac , \a_dinx[1]_cal1_u145_mac ,
       \a_dinx[1]_cal1_u146_mac , \a_dinx[1]_cal1_u147_mac , \a_dinx[1]_cal1_u148_mac ,
       \a_dinx[1]_cal1_u149_mac , \a_dinx[1]_coefcal1_u63_mac , \a_dinx[1]_coefcal1_u64_mac ,
       \a_dinx[1]_coefcal1_u64_mac_0_ , \a_dinx[2]_cal1_u137_mac , \a_dinx[2]_cal1_u138_mac ,
       \a_dinx[2]_cal1_u139_mac , \a_dinx[2]_cal1_u140_mac , \a_dinx[2]_cal1_u141_mac ,
       \a_dinx[2]_cal1_u142_mac , \a_dinx[2]_cal1_u143_mac , \a_dinx[2]_cal1_u144_mac ,
       \a_dinx[2]_cal1_u145_mac , \a_dinx[2]_cal1_u146_mac , \a_dinx[2]_cal1_u147_mac ,
       \a_dinx[2]_cal1_u148_mac , \a_dinx[2]_cal1_u149_mac , \a_dinx[2]_coefcal1_u63_mac ,
       \a_dinx[2]_coefcal1_u64_mac , \a_dinx[2]_coefcal1_u64_mac_0_ , \a_dinx[3]_cal1_u137_mac ,
       \a_dinx[3]_cal1_u138_mac , \a_dinx[3]_cal1_u139_mac , \a_dinx[3]_cal1_u140_mac ,
       \a_dinx[3]_cal1_u141_mac , \a_dinx[3]_cal1_u142_mac , \a_dinx[3]_cal1_u143_mac ,
       \a_dinx[3]_cal1_u144_mac , \a_dinx[3]_cal1_u145_mac , \a_dinx[3]_cal1_u146_mac ,
       \a_dinx[3]_cal1_u147_mac , \a_dinx[3]_cal1_u148_mac , \a_dinx[3]_cal1_u149_mac ,
       \a_dinx[3]_coefcal1_u63_mac , \a_dinx[3]_coefcal1_u64_mac , \a_dinx[3]_coefcal1_u64_mac_0_ ,
       \a_dinx[4]_cal1_u137_mac , \a_dinx[4]_cal1_u138_mac , \a_dinx[4]_cal1_u139_mac ,
       \a_dinx[4]_cal1_u140_mac , \a_dinx[4]_cal1_u141_mac , \a_dinx[4]_cal1_u142_mac ,
       \a_dinx[4]_cal1_u143_mac , \a_dinx[4]_cal1_u144_mac , \a_dinx[4]_cal1_u145_mac ,
       \a_dinx[4]_cal1_u146_mac , \a_dinx[4]_cal1_u147_mac , \a_dinx[4]_cal1_u148_mac ,
       \a_dinx[4]_cal1_u149_mac , \a_dinx[4]_coefcal1_u63_mac , \a_dinx[4]_coefcal1_u64_mac ,
       \a_dinx[4]_coefcal1_u64_mac_0_ , \a_dinx[5]_cal1_u137_mac , \a_dinx[5]_cal1_u138_mac ,
       \a_dinx[5]_cal1_u139_mac , \a_dinx[5]_cal1_u140_mac , \a_dinx[5]_cal1_u141_mac ,
       \a_dinx[5]_cal1_u142_mac , \a_dinx[5]_cal1_u143_mac , \a_dinx[5]_cal1_u144_mac ,
       \a_dinx[5]_cal1_u145_mac , \a_dinx[5]_cal1_u146_mac , \a_dinx[5]_cal1_u147_mac ,
       \a_dinx[5]_cal1_u148_mac , \a_dinx[5]_cal1_u149_mac , \a_dinx[5]_coefcal1_u63_mac ,
       \a_dinx[5]_coefcal1_u64_mac , \a_dinx[5]_coefcal1_u64_mac_0_ , \a_dinx[6]_cal1_u137_mac ,
       \a_dinx[6]_cal1_u138_mac , \a_dinx[6]_cal1_u139_mac , \a_dinx[6]_cal1_u140_mac ,
       \a_dinx[6]_cal1_u141_mac , \a_dinx[6]_cal1_u142_mac , \a_dinx[6]_cal1_u143_mac ,
       \a_dinx[6]_cal1_u144_mac , \a_dinx[6]_cal1_u145_mac , \a_dinx[6]_cal1_u146_mac ,
       \a_dinx[6]_cal1_u147_mac , \a_dinx[6]_cal1_u148_mac , \a_dinx[6]_cal1_u149_mac ,
       \a_dinx[6]_coefcal1_u63_mac , \a_dinx[6]_coefcal1_u64_mac , \a_dinx[6]_coefcal1_u64_mac_0_ ,
       \a_dinx[7]_cal1_u137_mac , \a_dinx[7]_cal1_u138_mac , \a_dinx[7]_cal1_u139_mac ,
       \a_dinx[7]_cal1_u140_mac , \a_dinx[7]_cal1_u141_mac , \a_dinx[7]_cal1_u142_mac ,
       \a_dinx[7]_cal1_u143_mac , \a_dinx[7]_cal1_u144_mac , \a_dinx[7]_cal1_u145_mac ,
       \a_dinx[7]_cal1_u146_mac , \a_dinx[7]_cal1_u147_mac , \a_dinx[7]_cal1_u148_mac ,
       \a_dinx[7]_cal1_u149_mac , \a_dinx[7]_coefcal1_u63_mac , \a_dinx[7]_coefcal1_u64_mac ,
       \a_dinx[7]_coefcal1_u64_mac_0_ , \a_dinx[8]_cal1_u137_mac , \a_dinx[8]_cal1_u138_mac ,
       \a_dinx[8]_cal1_u139_mac , \a_dinx[8]_cal1_u140_mac , \a_dinx[8]_cal1_u141_mac ,
       \a_dinx[8]_cal1_u142_mac , \a_dinx[8]_cal1_u143_mac , \a_dinx[8]_cal1_u144_mac ,
       \a_dinx[8]_cal1_u145_mac , \a_dinx[8]_cal1_u146_mac , \a_dinx[8]_cal1_u147_mac ,
       \a_dinx[8]_cal1_u148_mac , \a_dinx[8]_cal1_u149_mac , \a_dinx[8]_coefcal1_u63_mac ,
       \a_dinx[8]_coefcal1_u64_mac , \a_dinx[8]_coefcal1_u64_mac_0_ , \a_dinx[9]_cal1_u137_mac ,
       \a_dinx[9]_cal1_u138_mac , \a_dinx[9]_cal1_u139_mac , \a_dinx[9]_cal1_u140_mac ,
       \a_dinx[9]_cal1_u141_mac , \a_dinx[9]_cal1_u142_mac , \a_dinx[9]_cal1_u143_mac ,
       \a_dinx[9]_cal1_u144_mac , \a_dinx[9]_cal1_u145_mac , \a_dinx[9]_cal1_u146_mac ,
       \a_dinx[9]_cal1_u147_mac , \a_dinx[9]_cal1_u148_mac , \a_dinx[9]_cal1_u149_mac ,
       \a_dinx[9]_coefcal1_u63_mac , \a_dinx[9]_coefcal1_u64_mac , \a_dinx[9]_coefcal1_u64_mac_0_ ,
       a_dinxy_cen_cal1_u137_mac, a_dinxy_cen_cal1_u138_mac, a_dinxy_cen_cal1_u139_mac,
       a_dinxy_cen_cal1_u140_mac, a_dinxy_cen_cal1_u141_mac, a_dinxy_cen_cal1_u142_mac,
       a_dinxy_cen_cal1_u143_mac, a_dinxy_cen_cal1_u144_mac, a_dinxy_cen_cal1_u145_mac,
       a_dinxy_cen_cal1_u146_mac, a_dinxy_cen_cal1_u147_mac, a_dinxy_cen_cal1_u148_mac,
       a_dinxy_cen_cal1_u149_mac, a_dinxy_cen_coefcal1_u63_mac, a_dinxy_cen_coefcal1_u64_mac,
       a_dinxy_cen_coefcal1_u64_mac_0_, \a_diny[0]_cal1_u137_mac , \a_diny[0]_cal1_u138_mac ,
       \a_diny[0]_cal1_u139_mac , \a_diny[0]_cal1_u140_mac , \a_diny[0]_cal1_u141_mac ,
       \a_diny[0]_cal1_u142_mac , \a_diny[0]_cal1_u143_mac , \a_diny[0]_cal1_u144_mac ,
       \a_diny[0]_cal1_u145_mac , \a_diny[0]_cal1_u146_mac , \a_diny[0]_cal1_u147_mac ,
       \a_diny[0]_cal1_u148_mac , \a_diny[0]_cal1_u149_mac , \a_diny[0]_coefcal1_u63_mac ,
       \a_diny[0]_coefcal1_u64_mac , \a_diny[0]_coefcal1_u64_mac_0_ , \a_diny[1]_cal1_u137_mac ,
       \a_diny[1]_cal1_u138_mac , \a_diny[1]_cal1_u139_mac , \a_diny[1]_cal1_u140_mac ,
       \a_diny[1]_cal1_u141_mac , \a_diny[1]_cal1_u142_mac , \a_diny[1]_cal1_u143_mac ,
       \a_diny[1]_cal1_u144_mac , \a_diny[1]_cal1_u145_mac , \a_diny[1]_cal1_u146_mac ,
       \a_diny[1]_cal1_u147_mac , \a_diny[1]_cal1_u148_mac , \a_diny[1]_cal1_u149_mac ,
       \a_diny[1]_coefcal1_u63_mac , \a_diny[1]_coefcal1_u64_mac , \a_diny[1]_coefcal1_u64_mac_0_ ,
       \a_diny[2]_cal1_u137_mac , \a_diny[2]_cal1_u138_mac , \a_diny[2]_cal1_u139_mac ,
       \a_diny[2]_cal1_u140_mac , \a_diny[2]_cal1_u141_mac , \a_diny[2]_cal1_u142_mac ,
       \a_diny[2]_cal1_u143_mac , \a_diny[2]_cal1_u144_mac , \a_diny[2]_cal1_u145_mac ,
       \a_diny[2]_cal1_u146_mac , \a_diny[2]_cal1_u147_mac , \a_diny[2]_cal1_u148_mac ,
       \a_diny[2]_cal1_u149_mac , \a_diny[2]_coefcal1_u63_mac , \a_diny[2]_coefcal1_u64_mac ,
       \a_diny[2]_coefcal1_u64_mac_0_ , \a_diny[3]_cal1_u137_mac , \a_diny[3]_cal1_u138_mac ,
       \a_diny[3]_cal1_u139_mac , \a_diny[3]_cal1_u140_mac , \a_diny[3]_cal1_u141_mac ,
       \a_diny[3]_cal1_u142_mac , \a_diny[3]_cal1_u143_mac , \a_diny[3]_cal1_u144_mac ,
       \a_diny[3]_cal1_u145_mac , \a_diny[3]_cal1_u146_mac , \a_diny[3]_cal1_u147_mac ,
       \a_diny[3]_cal1_u148_mac , \a_diny[3]_cal1_u149_mac , \a_diny[3]_coefcal1_u63_mac ,
       \a_diny[3]_coefcal1_u64_mac , \a_diny[3]_coefcal1_u64_mac_0_ , \a_diny[4]_cal1_u137_mac ,
       \a_diny[4]_cal1_u138_mac , \a_diny[4]_cal1_u139_mac , \a_diny[4]_cal1_u140_mac ,
       \a_diny[4]_cal1_u141_mac , \a_diny[4]_cal1_u142_mac , \a_diny[4]_cal1_u143_mac ,
       \a_diny[4]_cal1_u144_mac , \a_diny[4]_cal1_u145_mac , \a_diny[4]_cal1_u146_mac ,
       \a_diny[4]_cal1_u147_mac , \a_diny[4]_cal1_u148_mac , \a_diny[4]_cal1_u149_mac ,
       \a_diny[4]_coefcal1_u63_mac , \a_diny[4]_coefcal1_u64_mac , \a_diny[4]_coefcal1_u64_mac_0_ ,
       \a_diny[5]_cal1_u137_mac , \a_diny[5]_cal1_u138_mac , \a_diny[5]_cal1_u139_mac ,
       \a_diny[5]_cal1_u140_mac , \a_diny[5]_cal1_u141_mac , \a_diny[5]_cal1_u142_mac ,
       \a_diny[5]_cal1_u143_mac , \a_diny[5]_cal1_u144_mac , \a_diny[5]_cal1_u145_mac ,
       \a_diny[5]_cal1_u146_mac , \a_diny[5]_cal1_u147_mac , \a_diny[5]_cal1_u148_mac ,
       \a_diny[5]_cal1_u149_mac , \a_diny[5]_coefcal1_u63_mac , \a_diny[5]_coefcal1_u64_mac ,
       \a_diny[5]_coefcal1_u64_mac_0_ , \a_diny[6]_cal1_u137_mac , \a_diny[6]_cal1_u138_mac ,
       \a_diny[6]_cal1_u139_mac , \a_diny[6]_cal1_u140_mac , \a_diny[6]_cal1_u141_mac ,
       \a_diny[6]_cal1_u142_mac , \a_diny[6]_cal1_u143_mac , \a_diny[6]_cal1_u144_mac ,
       \a_diny[6]_cal1_u145_mac , \a_diny[6]_cal1_u146_mac , \a_diny[6]_cal1_u147_mac ,
       \a_diny[6]_cal1_u148_mac , \a_diny[6]_cal1_u149_mac , \a_diny[6]_coefcal1_u63_mac ,
       \a_diny[6]_coefcal1_u64_mac , \a_diny[6]_coefcal1_u64_mac_0_ , \a_diny[7]_cal1_u137_mac ,
       \a_diny[7]_cal1_u138_mac , \a_diny[7]_cal1_u139_mac , \a_diny[7]_cal1_u140_mac ,
       \a_diny[7]_cal1_u141_mac , \a_diny[7]_cal1_u142_mac , \a_diny[7]_cal1_u143_mac ,
       \a_diny[7]_cal1_u144_mac , \a_diny[7]_cal1_u145_mac , \a_diny[7]_cal1_u146_mac ,
       \a_diny[7]_cal1_u147_mac , \a_diny[7]_cal1_u148_mac , \a_diny[7]_cal1_u149_mac ,
       \a_diny[7]_coefcal1_u63_mac , \a_diny[7]_coefcal1_u64_mac , \a_diny[7]_coefcal1_u64_mac_0_ ,
       \a_diny[8]_cal1_u137_mac , \a_diny[8]_cal1_u138_mac , \a_diny[8]_cal1_u139_mac ,
       \a_diny[8]_cal1_u140_mac , \a_diny[8]_cal1_u141_mac , \a_diny[8]_cal1_u142_mac ,
       \a_diny[8]_cal1_u143_mac , \a_diny[8]_cal1_u144_mac , \a_diny[8]_cal1_u145_mac ,
       \a_diny[8]_cal1_u146_mac , \a_diny[8]_cal1_u147_mac , \a_diny[8]_cal1_u148_mac ,
       \a_diny[8]_cal1_u149_mac , \a_diny[8]_coefcal1_u63_mac , \a_diny[8]_coefcal1_u64_mac ,
       \a_diny[8]_coefcal1_u64_mac_0_ , \a_diny[9]_cal1_u137_mac , \a_diny[9]_cal1_u138_mac ,
       \a_diny[9]_cal1_u139_mac , \a_diny[9]_cal1_u140_mac , \a_diny[9]_cal1_u141_mac ,
       \a_diny[9]_cal1_u142_mac , \a_diny[9]_cal1_u143_mac , \a_diny[9]_cal1_u144_mac ,
       \a_diny[9]_cal1_u145_mac , \a_diny[9]_cal1_u146_mac , \a_diny[9]_cal1_u147_mac ,
       \a_diny[9]_cal1_u148_mac , \a_diny[9]_cal1_u149_mac , \a_diny[9]_coefcal1_u63_mac ,
       \a_diny[9]_coefcal1_u64_mac , \a_diny[9]_coefcal1_u64_mac_0_ , a_dinz_cen_cal1_u137_mac,
       a_dinz_cen_cal1_u138_mac, a_dinz_cen_cal1_u139_mac, a_dinz_cen_cal1_u140_mac,
       a_dinz_cen_cal1_u141_mac, a_dinz_cen_cal1_u142_mac, a_dinz_cen_cal1_u143_mac,
       a_dinz_cen_cal1_u144_mac, a_dinz_cen_cal1_u145_mac, a_dinz_cen_cal1_u146_mac,
       a_dinz_cen_cal1_u147_mac, a_dinz_cen_cal1_u148_mac, a_dinz_cen_cal1_u149_mac,
       a_dinz_cen_coefcal1_u63_mac, a_dinz_cen_coefcal1_u64_mac, a_dinz_cen_coefcal1_u64_mac_0_,
       a_dinz_en_cal1_u137_mac, a_dinz_en_cal1_u138_mac, a_dinz_en_cal1_u139_mac,
       a_dinz_en_cal1_u140_mac, a_dinz_en_cal1_u141_mac, a_dinz_en_cal1_u142_mac,
       a_dinz_en_cal1_u143_mac, a_dinz_en_cal1_u144_mac, a_dinz_en_cal1_u145_mac,
       a_dinz_en_cal1_u146_mac, a_dinz_en_cal1_u147_mac, a_dinz_en_cal1_u148_mac,
       a_dinz_en_cal1_u149_mac, a_dinz_en_coefcal1_u63_mac, a_dinz_en_coefcal1_u64_mac,
       a_dinz_en_coefcal1_u64_mac_0_, a_in_sr_cal1_u137_mac, a_in_sr_cal1_u138_mac,
       a_in_sr_cal1_u139_mac, a_in_sr_cal1_u140_mac, a_in_sr_cal1_u141_mac, a_in_sr_cal1_u142_mac,
       a_in_sr_cal1_u143_mac, a_in_sr_cal1_u144_mac, a_in_sr_cal1_u145_mac, a_in_sr_cal1_u146_mac,
       a_in_sr_cal1_u147_mac, a_in_sr_cal1_u148_mac, a_in_sr_cal1_u149_mac, a_in_sr_coefcal1_u63_mac,
       a_in_sr_coefcal1_u64_mac, a_in_sr_coefcal1_u64_mac_0_;
    input  \a_mac_out[0]_coefcal1_u63_mac , \a_mac_out[0]_coefcal1_u64_mac ,
       \a_mac_out[0]_coefcal1_u64_mac_0_ , \a_mac_out[10]_cal1_u137_mac , \a_mac_out[10]_cal1_u138_mac ,
       \a_mac_out[10]_cal1_u139_mac , \a_mac_out[10]_cal1_u140_mac , \a_mac_out[10]_cal1_u141_mac ,
       \a_mac_out[10]_cal1_u142_mac , \a_mac_out[10]_cal1_u143_mac , \a_mac_out[10]_cal1_u144_mac ,
       \a_mac_out[10]_cal1_u145_mac , \a_mac_out[10]_cal1_u146_mac , \a_mac_out[10]_cal1_u147_mac ,
       \a_mac_out[10]_cal1_u148_mac , \a_mac_out[10]_cal1_u149_mac , \a_mac_out[10]_coefcal1_u63_mac ,
       \a_mac_out[10]_coefcal1_u64_mac , \a_mac_out[10]_coefcal1_u64_mac_0_ ,
       \a_mac_out[11]_cal1_u137_mac , \a_mac_out[11]_cal1_u138_mac , \a_mac_out[11]_cal1_u139_mac ,
       \a_mac_out[11]_cal1_u140_mac , \a_mac_out[11]_cal1_u141_mac , \a_mac_out[11]_cal1_u142_mac ,
       \a_mac_out[11]_cal1_u143_mac , \a_mac_out[11]_cal1_u144_mac , \a_mac_out[11]_cal1_u145_mac ,
       \a_mac_out[11]_cal1_u146_mac , \a_mac_out[11]_cal1_u147_mac , \a_mac_out[11]_cal1_u148_mac ,
       \a_mac_out[11]_cal1_u149_mac , \a_mac_out[11]_coefcal1_u63_mac , \a_mac_out[11]_coefcal1_u64_mac ,
       \a_mac_out[11]_coefcal1_u64_mac_0_ , \a_mac_out[12]_cal1_u138_mac , \a_mac_out[12]_cal1_u139_mac ,
       \a_mac_out[12]_cal1_u140_mac , \a_mac_out[12]_cal1_u141_mac , \a_mac_out[12]_cal1_u142_mac ,
       \a_mac_out[12]_cal1_u143_mac , \a_mac_out[12]_cal1_u144_mac , \a_mac_out[12]_cal1_u145_mac ,
       \a_mac_out[12]_cal1_u146_mac , \a_mac_out[12]_cal1_u147_mac , \a_mac_out[12]_cal1_u148_mac ,
       \a_mac_out[12]_cal1_u149_mac , \a_mac_out[12]_coefcal1_u63_mac , \a_mac_out[12]_coefcal1_u64_mac ,
       \a_mac_out[12]_coefcal1_u64_mac_0_ , \a_mac_out[13]_cal1_u138_mac , \a_mac_out[13]_cal1_u139_mac ,
       \a_mac_out[13]_cal1_u140_mac , \a_mac_out[13]_cal1_u141_mac , \a_mac_out[13]_cal1_u142_mac ,
       \a_mac_out[13]_cal1_u143_mac , \a_mac_out[13]_cal1_u144_mac , \a_mac_out[13]_cal1_u145_mac ,
       \a_mac_out[13]_cal1_u146_mac , \a_mac_out[13]_cal1_u147_mac , \a_mac_out[13]_cal1_u148_mac ,
       \a_mac_out[13]_cal1_u149_mac , \a_mac_out[13]_coefcal1_u63_mac , \a_mac_out[13]_coefcal1_u64_mac ,
       \a_mac_out[14]_coefcal1_u63_mac , \a_mac_out[14]_coefcal1_u64_mac , \a_mac_out[15]_coefcal1_u63_mac ,
       \a_mac_out[15]_coefcal1_u64_mac , \a_mac_out[16]_coefcal1_u63_mac , \a_mac_out[16]_coefcal1_u64_mac ,
       \a_mac_out[17]_coefcal1_u63_mac , \a_mac_out[17]_coefcal1_u64_mac , \a_mac_out[18]_coefcal1_u63_mac ,
       \a_mac_out[18]_coefcal1_u64_mac , \a_mac_out[19]_coefcal1_u63_mac , \a_mac_out[19]_coefcal1_u64_mac ,
       \a_mac_out[1]_coefcal1_u63_mac , \a_mac_out[1]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u64_mac_0_ ,
       \a_mac_out[20]_coefcal1_u64_mac , \a_mac_out[21]_coefcal1_u64_mac , \a_mac_out[22]_coefcal1_u64_mac ,
       \a_mac_out[23]_coefcal1_u64_mac , \a_mac_out[2]_coefcal1_u63_mac , \a_mac_out[2]_coefcal1_u64_mac ,
       \a_mac_out[2]_coefcal1_u64_mac_0_ , \a_mac_out[3]_coefcal1_u63_mac , \a_mac_out[3]_coefcal1_u64_mac ,
       \a_mac_out[3]_coefcal1_u64_mac_0_ , \a_mac_out[4]_coefcal1_u63_mac , \a_mac_out[4]_coefcal1_u64_mac ,
       \a_mac_out[4]_coefcal1_u64_mac_0_ , \a_mac_out[5]_coefcal1_u63_mac , \a_mac_out[5]_coefcal1_u64_mac ,
       \a_mac_out[5]_coefcal1_u64_mac_0_ , \a_mac_out[6]_cal1_u137_mac , \a_mac_out[6]_cal1_u138_mac ,
       \a_mac_out[6]_cal1_u139_mac , \a_mac_out[6]_cal1_u140_mac , \a_mac_out[6]_cal1_u141_mac ,
       \a_mac_out[6]_cal1_u142_mac , \a_mac_out[6]_cal1_u143_mac , \a_mac_out[6]_cal1_u144_mac ,
       \a_mac_out[6]_cal1_u145_mac , \a_mac_out[6]_cal1_u146_mac , \a_mac_out[6]_cal1_u147_mac ,
       \a_mac_out[6]_cal1_u148_mac , \a_mac_out[6]_cal1_u149_mac , \a_mac_out[6]_coefcal1_u63_mac ,
       \a_mac_out[6]_coefcal1_u64_mac , \a_mac_out[6]_coefcal1_u64_mac_0_ , \a_mac_out[7]_cal1_u137_mac ,
       \a_mac_out[7]_cal1_u138_mac , \a_mac_out[7]_cal1_u139_mac , \a_mac_out[7]_cal1_u140_mac ,
       \a_mac_out[7]_cal1_u141_mac , \a_mac_out[7]_cal1_u142_mac , \a_mac_out[7]_cal1_u143_mac ,
       \a_mac_out[7]_cal1_u144_mac , \a_mac_out[7]_cal1_u145_mac , \a_mac_out[7]_cal1_u146_mac ,
       \a_mac_out[7]_cal1_u147_mac , \a_mac_out[7]_cal1_u148_mac , \a_mac_out[7]_cal1_u149_mac ,
       \a_mac_out[7]_coefcal1_u63_mac , \a_mac_out[7]_coefcal1_u64_mac , \a_mac_out[7]_coefcal1_u64_mac_0_ ,
       \a_mac_out[8]_cal1_u137_mac , \a_mac_out[8]_cal1_u138_mac , \a_mac_out[8]_cal1_u139_mac ,
       \a_mac_out[8]_cal1_u140_mac , \a_mac_out[8]_cal1_u141_mac , \a_mac_out[8]_cal1_u142_mac ,
       \a_mac_out[8]_cal1_u143_mac , \a_mac_out[8]_cal1_u144_mac , \a_mac_out[8]_cal1_u145_mac ,
       \a_mac_out[8]_cal1_u146_mac , \a_mac_out[8]_cal1_u147_mac , \a_mac_out[8]_cal1_u148_mac ,
       \a_mac_out[8]_cal1_u149_mac , \a_mac_out[8]_coefcal1_u63_mac , \a_mac_out[8]_coefcal1_u64_mac ,
       \a_mac_out[8]_coefcal1_u64_mac_0_ , \a_mac_out[9]_cal1_u137_mac , \a_mac_out[9]_cal1_u138_mac ,
       \a_mac_out[9]_cal1_u139_mac , \a_mac_out[9]_cal1_u140_mac , \a_mac_out[9]_cal1_u141_mac ,
       \a_mac_out[9]_cal1_u142_mac , \a_mac_out[9]_cal1_u143_mac , \a_mac_out[9]_cal1_u144_mac ,
       \a_mac_out[9]_cal1_u145_mac , \a_mac_out[9]_cal1_u146_mac , \a_mac_out[9]_cal1_u147_mac ,
       \a_mac_out[9]_cal1_u148_mac , \a_mac_out[9]_cal1_u149_mac , \a_mac_out[9]_coefcal1_u63_mac ,
       \a_mac_out[9]_coefcal1_u64_mac , \a_mac_out[9]_coefcal1_u64_mac_0_ ;
    output a_mac_out_cen_cal1_u137_mac, a_mac_out_cen_cal1_u138_mac, a_mac_out_cen_cal1_u139_mac,
       a_mac_out_cen_cal1_u140_mac, a_mac_out_cen_cal1_u141_mac, a_mac_out_cen_cal1_u142_mac,
       a_mac_out_cen_cal1_u143_mac, a_mac_out_cen_cal1_u144_mac, a_mac_out_cen_cal1_u145_mac,
       a_mac_out_cen_cal1_u146_mac, a_mac_out_cen_cal1_u147_mac, a_mac_out_cen_cal1_u148_mac,
       a_mac_out_cen_cal1_u149_mac, a_mac_out_cen_coefcal1_u63_mac, a_mac_out_cen_coefcal1_u64_mac,
       a_mac_out_cen_coefcal1_u64_mac_0_, a_out_sr_cal1_u137_mac, a_out_sr_cal1_u138_mac,
       a_out_sr_cal1_u139_mac, a_out_sr_cal1_u140_mac, a_out_sr_cal1_u141_mac,
       a_out_sr_cal1_u142_mac, a_out_sr_cal1_u143_mac, a_out_sr_cal1_u144_mac,
       a_out_sr_cal1_u145_mac, a_out_sr_cal1_u146_mac, a_out_sr_cal1_u147_mac,
       a_out_sr_cal1_u148_mac, a_out_sr_cal1_u149_mac, a_out_sr_coefcal1_u63_mac,
       a_out_sr_coefcal1_u64_mac, a_out_sr_coefcal1_u64_mac_0_, a_sload_cal1_u137_mac,
       a_sload_cal1_u138_mac, a_sload_cal1_u139_mac, a_sload_cal1_u140_mac, a_sload_cal1_u141_mac,
       a_sload_cal1_u142_mac, a_sload_cal1_u143_mac, a_sload_cal1_u144_mac, a_sload_cal1_u145_mac,
       a_sload_cal1_u146_mac, a_sload_cal1_u147_mac, a_sload_cal1_u148_mac, a_sload_cal1_u149_mac,
       a_sload_coefcal1_u63_mac, a_sload_coefcal1_u64_mac, a_sload_coefcal1_u64_mac_0_,
       b_acc_en_coefcal1_u64_mac, b_acc_en_coefcal1_u64_mac_0_, \b_dinx[0]_coefcal1_u64_mac ,
       \b_dinx[0]_coefcal1_u64_mac_0_ , \b_dinx[10]_coefcal1_u64_mac , \b_dinx[10]_coefcal1_u64_mac_0_ ,
       \b_dinx[11]_coefcal1_u64_mac , \b_dinx[11]_coefcal1_u64_mac_0_ , \b_dinx[12]_coefcal1_u64_mac ,
       \b_dinx[12]_coefcal1_u64_mac_0_ , \b_dinx[13]_coefcal1_u64_mac , \b_dinx[13]_coefcal1_u64_mac_0_ ,
       \b_dinx[1]_coefcal1_u64_mac , \b_dinx[1]_coefcal1_u64_mac_0_ , \b_dinx[2]_coefcal1_u64_mac ,
       \b_dinx[2]_coefcal1_u64_mac_0_ , \b_dinx[3]_coefcal1_u64_mac , \b_dinx[3]_coefcal1_u64_mac_0_ ,
       \b_dinx[4]_coefcal1_u64_mac , \b_dinx[4]_coefcal1_u64_mac_0_ , \b_dinx[5]_coefcal1_u64_mac ,
       \b_dinx[5]_coefcal1_u64_mac_0_ , \b_dinx[6]_coefcal1_u64_mac , \b_dinx[6]_coefcal1_u64_mac_0_ ,
       \b_dinx[7]_coefcal1_u64_mac , \b_dinx[7]_coefcal1_u64_mac_0_ , \b_dinx[8]_coefcal1_u64_mac ,
       \b_dinx[8]_coefcal1_u64_mac_0_ , \b_dinx[9]_coefcal1_u64_mac , \b_dinx[9]_coefcal1_u64_mac_0_ ,
       b_dinxy_cen_coefcal1_u64_mac, b_dinxy_cen_coefcal1_u64_mac_0_, \b_diny[0]_coefcal1_u64_mac ,
       \b_diny[0]_coefcal1_u64_mac_0_ , \b_diny[1]_coefcal1_u64_mac , \b_diny[1]_coefcal1_u64_mac_0_ ,
       \b_diny[2]_coefcal1_u64_mac , \b_diny[2]_coefcal1_u64_mac_0_ , \b_diny[3]_coefcal1_u64_mac ,
       \b_diny[3]_coefcal1_u64_mac_0_ , \b_diny[4]_coefcal1_u64_mac , \b_diny[4]_coefcal1_u64_mac_0_ ,
       \b_diny[5]_coefcal1_u64_mac , \b_diny[5]_coefcal1_u64_mac_0_ , \b_diny[6]_coefcal1_u64_mac ,
       \b_diny[6]_coefcal1_u64_mac_0_ , \b_diny[7]_coefcal1_u64_mac , \b_diny[7]_coefcal1_u64_mac_0_ ,
       \b_diny[8]_coefcal1_u64_mac , \b_diny[8]_coefcal1_u64_mac_0_ , \b_diny[9]_coefcal1_u64_mac ,
       \b_diny[9]_coefcal1_u64_mac_0_ , b_dinz_cen_coefcal1_u64_mac, b_dinz_cen_coefcal1_u64_mac_0_,
       b_dinz_en_coefcal1_u64_mac, b_dinz_en_coefcal1_u64_mac_0_, b_in_sr_coefcal1_u64_mac,
       b_in_sr_coefcal1_u64_mac_0_;
    input  \b_mac_out[0]_coefcal1_u64_mac , \b_mac_out[1]_coefcal1_u64_mac ,
       \b_mac_out[2]_coefcal1_u64_mac , \b_mac_out[3]_coefcal1_u64_mac , \b_mac_out[4]_coefcal1_u64_mac ;
    output b_mac_out_cen_coefcal1_u64_mac, b_mac_out_cen_coefcal1_u64_mac_0_,
       b_out_sr_coefcal1_u64_mac, b_out_sr_coefcal1_u64_mac_0_, b_sload_coefcal1_u64_mac,
       b_sload_coefcal1_u64_mac_0_, \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_1 , c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_0A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_0B_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_0B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_1A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_1B_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_1B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2A_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_2A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_2B_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_2B_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3A_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_3A_u_emb18k_1, c1r1_clka_fifo1_ram_inst_3B_u_emb18k_0,
       c1r1_clka_fifo1_ram_inst_3B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_1, c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_0,
       c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_1, \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_1 , \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    input  \c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r1_q[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r1_q[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    output c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_1,
       c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_0, c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_0, c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_0A_u_emb18k_0, c1r2_clka_fifo1_ram_inst_0A_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_0B_u_emb18k_0, c1r2_clka_fifo1_ram_inst_0B_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_1A_u_emb18k_0, c1r2_clka_fifo1_ram_inst_1A_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_1B_u_emb18k_0, c1r2_clka_fifo1_ram_inst_1B_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_2A_u_emb18k_0, c1r2_clka_fifo1_ram_inst_2A_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_2B_u_emb18k_0, c1r2_clka_fifo1_ram_inst_2B_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_3A_u_emb18k_0, c1r2_clka_fifo1_ram_inst_3A_u_emb18k_1,
       c1r2_clka_fifo1_ram_inst_3B_u_emb18k_0, c1r2_clka_fifo1_ram_inst_3B_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_0, c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_1,
       \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    input  \c1r2_q[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r2_q[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r2_q[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r2_q[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r2_q[9]_fifo1_ram_inst_3B_u_emb18k_0 ;
    output c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_1,
       c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_0, c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_0, c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_0A_u_emb18k_0, c1r3_clka_fifo1_ram_inst_0A_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_0B_u_emb18k_0, c1r3_clka_fifo1_ram_inst_0B_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_1A_u_emb18k_0, c1r3_clka_fifo1_ram_inst_1A_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_1B_u_emb18k_0, c1r3_clka_fifo1_ram_inst_1B_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_2A_u_emb18k_0, c1r3_clka_fifo1_ram_inst_2A_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_2B_u_emb18k_0, c1r3_clka_fifo1_ram_inst_2B_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_3A_u_emb18k_0, c1r3_clka_fifo1_ram_inst_3A_u_emb18k_1,
       c1r3_clka_fifo1_ram_inst_3B_u_emb18k_0, c1r3_clka_fifo1_ram_inst_3B_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_0, c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_1,
       \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    input  \c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r3_q[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r3_q[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    output c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_1,
       c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_0, c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_0, c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_0A_u_emb18k_0, c1r4_clka_fifo1_ram_inst_0A_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_0B_u_emb18k_0, c1r4_clka_fifo1_ram_inst_0B_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_1A_u_emb18k_0, c1r4_clka_fifo1_ram_inst_1A_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_1B_u_emb18k_0, c1r4_clka_fifo1_ram_inst_1B_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_2A_u_emb18k_0, c1r4_clka_fifo1_ram_inst_2A_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_2B_u_emb18k_0, c1r4_clka_fifo1_ram_inst_2B_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_3A_u_emb18k_0, c1r4_clka_fifo1_ram_inst_3A_u_emb18k_1,
       c1r4_clka_fifo1_ram_inst_3B_u_emb18k_0, c1r4_clka_fifo1_ram_inst_3B_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_0, c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_1,
       \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_0 , \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_1 ;
    input  \c1r4_q[0]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[0]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[0]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[0]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[10]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[10]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[10]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[10]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[11]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[11]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[11]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[11]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[12]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[12]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[12]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[12]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[1]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[1]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[1]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[1]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[2]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[2]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[2]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[2]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[3]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[3]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[3]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[3]_fifo1_ram_inst_3B_u_emb18k_0 ,
       \c1r4_q[9]_fifo1_ram_inst_0A_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ,
       \c1r4_q[9]_fifo1_ram_inst_1A_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ,
       \c1r4_q[9]_fifo1_ram_inst_3A_u_emb18k_0 , \c1r4_q[9]_fifo1_ram_inst_3B_u_emb18k_0 ;
    output c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_1,
       c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_0, c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_1,
       c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_0, c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_1,
       cea_fifo1_ram_inst_0A_u_emb18k_0, cea_fifo1_ram_inst_0A_u_emb18k_1, cea_fifo1_ram_inst_0B_u_emb18k_0,
       cea_fifo1_ram_inst_0B_u_emb18k_1, cea_fifo1_ram_inst_1A_u_emb18k_0, cea_fifo1_ram_inst_1A_u_emb18k_1,
       cea_fifo1_ram_inst_1B_u_emb18k_0, cea_fifo1_ram_inst_1B_u_emb18k_1, cea_fifo1_ram_inst_2A_u_emb18k_0,
       cea_fifo1_ram_inst_2A_u_emb18k_1, cea_fifo1_ram_inst_2B_u_emb18k_0, cea_fifo1_ram_inst_2B_u_emb18k_1,
       cea_fifo1_ram_inst_3A_u_emb18k_0, cea_fifo1_ram_inst_3A_u_emb18k_1, cea_fifo1_ram_inst_3B_u_emb18k_0,
       cea_fifo1_ram_inst_3B_u_emb18k_1, ceb_fifo1_ram_inst_0A_u_emb18k_0, ceb_fifo1_ram_inst_0A_u_emb18k_1,
       ceb_fifo1_ram_inst_0B_u_emb18k_0, ceb_fifo1_ram_inst_0B_u_emb18k_1, ceb_fifo1_ram_inst_1A_u_emb18k_0,
       ceb_fifo1_ram_inst_1A_u_emb18k_1, ceb_fifo1_ram_inst_1B_u_emb18k_0, ceb_fifo1_ram_inst_1B_u_emb18k_1,
       ceb_fifo1_ram_inst_2A_u_emb18k_0, ceb_fifo1_ram_inst_2A_u_emb18k_1, ceb_fifo1_ram_inst_2B_u_emb18k_0,
       ceb_fifo1_ram_inst_2B_u_emb18k_1, ceb_fifo1_ram_inst_3A_u_emb18k_0, ceb_fifo1_ram_inst_3A_u_emb18k_1,
       ceb_fifo1_ram_inst_3B_u_emb18k_0, ceb_fifo1_ram_inst_3B_u_emb18k_1;
    input  clka, clkb;
    input  [23:0] dIn;
    input  dInEn;
    output [23:0] dOut;
    output dOutEn;
    input  en;
    output \haa[0]_fifo1_ram_inst_0A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_0B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_1B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_2A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_2B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_3A_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \haa[0]_fifo1_ram_inst_3B_u_emb18k_0 , \haa[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_0A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_0B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_1A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_1B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_2A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_2B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_3A_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \haa[1]_fifo1_ram_inst_3B_u_emb18k_0 , \haa[1]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_0A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_0B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_1A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_1B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_2A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_2B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_3A_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \hab[0]_fifo1_ram_inst_3B_u_emb18k_0 , \hab[0]_fifo1_ram_inst_3B_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_0A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0A_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_0B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_0B_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_1A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1A_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_1B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_1B_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_2A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2A_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_2B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_2B_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_3A_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3A_u_emb18k_1 ,
       \hab[1]_fifo1_ram_inst_3B_u_emb18k_0 , \hab[1]_fifo1_ram_inst_3B_u_emb18k_1 ;
    input  iHsyn, iVsyn;
    input  [10:0] inXRes;
    input  [10:0] inYRes;
    input  [11:0] outXRes;
    input  [11:0] outYRes;
    input  rst;
    output u5018_OUT;
    input  u5502_I1, u5502_I1_5_, u5502_IN, u5859_I1;
    output u8205_O, u8205_O_1_, u8205_O_2_, u8218_Y, u8224_O, u8224_O_4_, u8230_O,
       u8231_O;
    input  u8245_D0, u8245_I0, u8245_I0_0_, u8245_I0_3_, u8245_IN;
    output wea_fifo1_ram_inst_0A_u_emb18k_0, wea_fifo1_ram_inst_0A_u_emb18k_1,
       wea_fifo1_ram_inst_0B_u_emb18k_0, wea_fifo1_ram_inst_0B_u_emb18k_1, wea_fifo1_ram_inst_1A_u_emb18k_0,
       wea_fifo1_ram_inst_1A_u_emb18k_1, wea_fifo1_ram_inst_1B_u_emb18k_0, wea_fifo1_ram_inst_1B_u_emb18k_1,
       wea_fifo1_ram_inst_2A_u_emb18k_0, wea_fifo1_ram_inst_2A_u_emb18k_1, wea_fifo1_ram_inst_2B_u_emb18k_0,
       wea_fifo1_ram_inst_2B_u_emb18k_1, wea_fifo1_ram_inst_3A_u_emb18k_0, wea_fifo1_ram_inst_3A_u_emb18k_1,
       wea_fifo1_ram_inst_3B_u_emb18k_0, wea_fifo1_ram_inst_3B_u_emb18k_1, web_fifo1_ram_inst_0A_u_emb18k_0,
       web_fifo1_ram_inst_0A_u_emb18k_1, web_fifo1_ram_inst_0B_u_emb18k_0, web_fifo1_ram_inst_0B_u_emb18k_1,
       web_fifo1_ram_inst_1A_u_emb18k_0, web_fifo1_ram_inst_1A_u_emb18k_1, web_fifo1_ram_inst_1B_u_emb18k_0,
       web_fifo1_ram_inst_1B_u_emb18k_1, web_fifo1_ram_inst_2A_u_emb18k_0, web_fifo1_ram_inst_2A_u_emb18k_1,
       web_fifo1_ram_inst_2B_u_emb18k_0, web_fifo1_ram_inst_2B_u_emb18k_1, web_fifo1_ram_inst_3A_u_emb18k_0,
       web_fifo1_ram_inst_3A_u_emb18k_1, web_fifo1_ram_inst_3B_u_emb18k_0, web_fifo1_ram_inst_3B_u_emb18k_1;
    input  [10:0] xBgn;
    input  [10:0] xEnd;
    input  [10:0] yBgn;
    input  [10:0] yEnd;
    wire   HS_2079_net, \cal1_VSNormal__reg|Q_net , \cal1_enforceJmp__reg|Q_net ,
       \cal1_jmp1Normal__reg|Q_net , \cal1_jmp2Normal__reg|Q_net , \cal1_ramRdAddr__reg[0]|Q_net ,
       \cal1_ramRdAddr__reg[10]|Q_net , \cal1_ramRdAddr__reg[1]|Q_net , \cal1_ramRdAddr__reg[2]|Q_net ,
       \cal1_ramRdAddr__reg[3]|Q_net , \cal1_ramRdAddr__reg[4]|Q_net , \cal1_ramRdAddr__reg[5]|Q_net ,
       \cal1_ramRdAddr__reg[6]|Q_net , \cal1_ramRdAddr__reg[7]|Q_net , \cal1_ramRdAddr__reg[8]|Q_net ,
       \cal1_ramRdAddr__reg[9]|Q_net , \cal1_u127_XORCI_0|SUM_net , \cal1_u127_XORCI_10|SUM_net ,
       \cal1_u127_XORCI_11|SUM_net , \cal1_u127_XORCI_12|SUM_net , \cal1_u127_XORCI_13|SUM_net ,
       \cal1_u127_XORCI_14|SUM_net , \cal1_u127_XORCI_15|SUM_net , \cal1_u127_XORCI_16|SUM_net ,
       \cal1_u127_XORCI_1|SUM_net , \cal1_u127_XORCI_2|SUM_net , \cal1_u127_XORCI_3|SUM_net ,
       \cal1_u127_XORCI_4|SUM_net , \cal1_u127_XORCI_5|SUM_net , \cal1_u127_XORCI_6|SUM_net ,
       \cal1_u127_XORCI_7|SUM_net , \cal1_u127_XORCI_8|SUM_net , \cal1_u127_XORCI_9|SUM_net ,
       \cal1_u128_XORCI_0|SUM_net , \cal1_u128_XORCI_10|SUM_net , \cal1_u128_XORCI_11|SUM_net ,
       \cal1_u128_XORCI_12|SUM_net , \cal1_u128_XORCI_13|SUM_net , \cal1_u128_XORCI_14|SUM_net ,
       \cal1_u128_XORCI_15|SUM_net , \cal1_u128_XORCI_16|SUM_net , \cal1_u128_XORCI_1|SUM_net ,
       \cal1_u128_XORCI_2|SUM_net , \cal1_u128_XORCI_3|SUM_net , \cal1_u128_XORCI_4|SUM_net ,
       \cal1_u128_XORCI_5|SUM_net , \cal1_u128_XORCI_6|SUM_net , \cal1_u128_XORCI_7|SUM_net ,
       \cal1_u128_XORCI_8|SUM_net , \cal1_u128_XORCI_9|SUM_net , \cal1_u129_XORCI_0|SUM_net ,
       \cal1_u129_XORCI_10|SUM_net , \cal1_u129_XORCI_1|SUM_net , \cal1_u129_XORCI_2|SUM_net ,
       \cal1_u129_XORCI_3|SUM_net , \cal1_u129_XORCI_4|SUM_net , \cal1_u129_XORCI_5|SUM_net ,
       \cal1_u129_XORCI_6|SUM_net , \cal1_u129_XORCI_7|SUM_net , \cal1_u129_XORCI_8|SUM_net ,
       \cal1_u129_XORCI_9|SUM_net , \cal1_u130_XORCI_0|SUM_net , \cal1_u130_XORCI_10|SUM_net ,
       \cal1_u130_XORCI_1|SUM_net , \cal1_u130_XORCI_2|SUM_net , \cal1_u130_XORCI_3|SUM_net ,
       \cal1_u130_XORCI_4|SUM_net , \cal1_u130_XORCI_5|SUM_net , \cal1_u130_XORCI_6|SUM_net ,
       \cal1_u130_XORCI_7|SUM_net , \cal1_u130_XORCI_8|SUM_net , \cal1_u130_XORCI_9|SUM_net ,
       \cal1_u131_XORCI_0|SUM_net , \cal1_u131_XORCI_10|SUM_net , \cal1_u131_XORCI_1|SUM_net ,
       \cal1_u131_XORCI_2|SUM_net , \cal1_u131_XORCI_3|SUM_net , \cal1_u131_XORCI_4|SUM_net ,
       \cal1_u131_XORCI_5|SUM_net , \cal1_u131_XORCI_6|SUM_net , \cal1_u131_XORCI_7|SUM_net ,
       \cal1_u131_XORCI_8|SUM_net , \cal1_u131_XORCI_9|SUM_net , \cal1_u132_XORCI_0|SUM_net ,
       \cal1_u132_XORCI_10|SUM_net , \cal1_u132_XORCI_1|SUM_net , \cal1_u132_XORCI_2|SUM_net ,
       \cal1_u132_XORCI_3|SUM_net , \cal1_u132_XORCI_4|SUM_net , \cal1_u132_XORCI_5|SUM_net ,
       \cal1_u132_XORCI_6|SUM_net , \cal1_u132_XORCI_7|SUM_net , \cal1_u132_XORCI_8|SUM_net ,
       \cal1_u132_XORCI_9|SUM_net , \cal1_u133_XORCI_0|SUM_net , \cal1_u133_XORCI_1|SUM_net ,
       \cal1_u133_XORCI_2|SUM_net , \cal1_u133_XORCI_3|SUM_net , \cal1_u133_XORCI_4|SUM_net ,
       \cal1_u133_XORCI_5|SUM_net , \cal1_u133_XORCI_6|SUM_net , \cal1_u134_SUM_XORCI_0_10_|SUM_net ,
       \cal1_u134_SUM_XORCI_0_13_|SUM_net , \cal1_u134_SUM_XORCI_0_16_|SUM_net ,
       \cal1_u134_SUM_XORCI_0_19_|SUM_net , \cal1_u134_SUM_XORCI_0_1_|SUM_net ,
       \cal1_u134_SUM_XORCI_0_4_|SUM_net , \cal1_u134_SUM_XORCI_0_7_|SUM_net ,
       \cal1_u134_SUM_XORCI_0|SUM_net , \cal1_u134_SUM_XORCI_1_22_|SUM_net ,
       \cal1_u134_SUM_XORCI_1_25_|SUM_net , \cal1_u134_SUM_XORCI_1_28_|SUM_net ,
       \cal1_u134_SUM_XORCI_1_31_|SUM_net , \cal1_u134_SUM_XORCI_1_34_|SUM_net ,
       \cal1_u134_SUM_XORCI_1_37_|SUM_net , \cal1_u134_SUM_XORCI_1_40_|SUM_net ,
       \cal1_u134_SUM_XORCI_1|SUM_net , \cal1_u134_XORCI_SHIFT_0|SUM_net , \cal1_u134_XORCI_SHIFT_1|SUM_net ,
       \cal1_u135_SUM_XORCI_0_67_|SUM_net , \cal1_u135_SUM_XORCI_0_70_|SUM_net ,
       \cal1_u135_SUM_XORCI_0_73_|SUM_net , \cal1_u135_SUM_XORCI_0_76_|SUM_net ,
       \cal1_u135_SUM_XORCI_0_79_|SUM_net , \cal1_u135_SUM_XORCI_0_82_|SUM_net ,
       \cal1_u135_SUM_XORCI_0_85_|SUM_net , \cal1_u135_SUM_XORCI_0|SUM_net ,
       \cal1_u135_SUM_XORCI_1_100_|SUM_net , \cal1_u135_SUM_XORCI_1_103_|SUM_net ,
       \cal1_u135_SUM_XORCI_1_106_|SUM_net , \cal1_u135_SUM_XORCI_1_88_|SUM_net ,
       \cal1_u135_SUM_XORCI_1_91_|SUM_net , \cal1_u135_SUM_XORCI_1_94_|SUM_net ,
       \cal1_u135_SUM_XORCI_1_97_|SUM_net , \cal1_u135_SUM_XORCI_1|SUM_net ,
       \cal1_u135_XORCI_SHIFT_0|SUM_net , \cal1_u135_XORCI_SHIFT_1|SUM_net ,
       \cal1_u136_SUM_XORCI_0_133_|SUM_net , \cal1_u136_SUM_XORCI_0_136_|SUM_net ,
       \cal1_u136_SUM_XORCI_0_139_|SUM_net , \cal1_u136_SUM_XORCI_0_142_|SUM_net ,
       \cal1_u136_SUM_XORCI_0_145_|SUM_net , \cal1_u136_SUM_XORCI_0_148_|SUM_net ,
       \cal1_u136_SUM_XORCI_0_151_|SUM_net , \cal1_u136_SUM_XORCI_0|SUM_net ,
       \cal1_u136_SUM_XORCI_1_154_|SUM_net , \cal1_u136_SUM_XORCI_1_157_|SUM_net ,
       \cal1_u136_SUM_XORCI_1_160_|SUM_net , \cal1_u136_SUM_XORCI_1_163_|SUM_net ,
       \cal1_u136_SUM_XORCI_1_166_|SUM_net , \cal1_u136_SUM_XORCI_1_169_|SUM_net ,
       \cal1_u136_SUM_XORCI_1_172_|SUM_net , \cal1_u136_SUM_XORCI_1|SUM_net ,
       \cal1_u136_XORCI_SHIFT_0|SUM_net , \cal1_u136_XORCI_SHIFT_1|SUM_net ,
       \cal1_u54_XORCI_0|SUM_net , \cal1_u54_XORCI_1|SUM_net , \cal1_u54_XORCI_2|SUM_net ,
       \cal1_u54_XORCI_3|SUM_net , \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_5|SUM_net ,
       \cal1_u54_XORCI_6|SUM_net , \cal1_u55_XORCI_0|SUM_net , \cal1_u55_XORCI_1|SUM_net ,
       \cal1_u55_XORCI_2|SUM_net , \cal1_u55_XORCI_3|SUM_net , \cal1_u55_XORCI_4|SUM_net ,
       \cal1_u55_XORCI_5|SUM_net , \cal1_u55_XORCI_6|SUM_net , \cal1_u57_XORCI_11|SUM_net ,
       \cal1_u59_XORCI_11|SUM_net , \cal1_u61_XORCI_11|SUM_net , \cal1_u63_XORCI_11|SUM_net ,
       \cal1_uPreF__reg[0]|Q_net , \cal1_uPreF__reg[1]|Q_net , \cal1_uPreF__reg[2]|Q_net ,
       \cal1_uPreF__reg[3]|Q_net , \cal1_uPreF__reg[4]|Q_net , \cal1_uPreF__reg[5]|Q_net ,
       \cal1_u__reg[0]|Q_net , \cal1_u__reg[10]|Q_net , \cal1_u__reg[11]|Q_net ,
       \cal1_u__reg[12]|Q_net , \cal1_u__reg[13]|Q_net , \cal1_u__reg[14]|Q_net ,
       \cal1_u__reg[15]|Q_net , \cal1_u__reg[16]|Q_net , \cal1_u__reg[1]|Q_net ,
       \cal1_u__reg[2]|Q_net , \cal1_u__reg[3]|Q_net , \cal1_u__reg[4]|Q_net ,
       \cal1_u__reg[5]|Q_net , \cal1_u__reg[6]|Q_net , \cal1_u__reg[7]|Q_net ,
       \cal1_u__reg[8]|Q_net , \cal1_u__reg[9]|Q_net , \cal1_v__reg[0]|Q_net ,
       \cal1_v__reg[10]|Q_net , \cal1_v__reg[11]|Q_net , \cal1_v__reg[12]|Q_net ,
       \cal1_v__reg[13]|Q_net , \cal1_v__reg[14]|Q_net , \cal1_v__reg[15]|Q_net ,
       \cal1_v__reg[16]|Q_net , \cal1_v__reg[1]|Q_net , \cal1_v__reg[2]|Q_net ,
       \cal1_v__reg[3]|Q_net , \cal1_v__reg[4]|Q_net , \cal1_v__reg[5]|Q_net ,
       \cal1_v__reg[6]|Q_net , \cal1_v__reg[7]|Q_net , \cal1_v__reg[8]|Q_net ,
       \cal1_v__reg[9]|Q_net , \cal1_xAddress__reg[0]|Q_net , \cal1_xAddress__reg[10]|Q_net ,
       \cal1_xAddress__reg[1]|Q_net , \cal1_xAddress__reg[2]|Q_net , \cal1_xAddress__reg[3]|Q_net ,
       \cal1_xAddress__reg[4]|Q_net , \cal1_xAddress__reg[5]|Q_net , \cal1_xAddress__reg[6]|Q_net ,
       \cal1_xAddress__reg[7]|Q_net , \cal1_xAddress__reg[8]|Q_net , \cal1_xAddress__reg[9]|Q_net ,
       \cal1_yAddress__reg[0]|Q_net , \cal1_yAddress__reg[10]|Q_net , \cal1_yAddress__reg[1]|Q_net ,
       \cal1_yAddress__reg[2]|Q_net , \cal1_yAddress__reg[3]|Q_net , \cal1_yAddress__reg[4]|Q_net ,
       \cal1_yAddress__reg[5]|Q_net , \cal1_yAddress__reg[6]|Q_net , \cal1_yAddress__reg[7]|Q_net ,
       \cal1_yAddress__reg[8]|Q_net , \cal1_yAddress__reg[9]|Q_net , \coefcal1_divide_inst1_u102_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_10|SUM_net , \coefcal1_divide_inst1_u102_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_12|SUM_net , \coefcal1_divide_inst1_u102_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_14|SUM_net , \coefcal1_divide_inst1_u102_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_1|SUM_net , \coefcal1_divide_inst1_u102_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_3|SUM_net , \coefcal1_divide_inst1_u102_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_5|SUM_net , \coefcal1_divide_inst1_u102_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_7|SUM_net , \coefcal1_divide_inst1_u102_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u102_XORCI_9|SUM_net , \coefcal1_divide_inst1_u103_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_10|SUM_net , \coefcal1_divide_inst1_u103_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_12|SUM_net , \coefcal1_divide_inst1_u103_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_14|SUM_net , \coefcal1_divide_inst1_u103_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_1|SUM_net , \coefcal1_divide_inst1_u103_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_3|SUM_net , \coefcal1_divide_inst1_u103_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_5|SUM_net , \coefcal1_divide_inst1_u103_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_7|SUM_net , \coefcal1_divide_inst1_u103_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u103_XORCI_9|SUM_net , \coefcal1_divide_inst1_u104_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_10|SUM_net , \coefcal1_divide_inst1_u104_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_12|SUM_net , \coefcal1_divide_inst1_u104_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_14|SUM_net , \coefcal1_divide_inst1_u104_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_1|SUM_net , \coefcal1_divide_inst1_u104_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_3|SUM_net , \coefcal1_divide_inst1_u104_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_5|SUM_net , \coefcal1_divide_inst1_u104_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_7|SUM_net , \coefcal1_divide_inst1_u104_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u104_XORCI_9|SUM_net , \coefcal1_divide_inst1_u105_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_10|SUM_net , \coefcal1_divide_inst1_u105_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_12|SUM_net , \coefcal1_divide_inst1_u105_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_14|SUM_net , \coefcal1_divide_inst1_u105_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_1|SUM_net , \coefcal1_divide_inst1_u105_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_3|SUM_net , \coefcal1_divide_inst1_u105_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_5|SUM_net , \coefcal1_divide_inst1_u105_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_7|SUM_net , \coefcal1_divide_inst1_u105_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u105_XORCI_9|SUM_net , \coefcal1_divide_inst1_u106_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_10|SUM_net , \coefcal1_divide_inst1_u106_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_12|SUM_net , \coefcal1_divide_inst1_u106_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_14|SUM_net , \coefcal1_divide_inst1_u106_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_1|SUM_net , \coefcal1_divide_inst1_u106_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_3|SUM_net , \coefcal1_divide_inst1_u106_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_5|SUM_net , \coefcal1_divide_inst1_u106_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_7|SUM_net , \coefcal1_divide_inst1_u106_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u106_XORCI_9|SUM_net , \coefcal1_divide_inst1_u107_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_10|SUM_net , \coefcal1_divide_inst1_u107_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_12|SUM_net , \coefcal1_divide_inst1_u107_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_14|SUM_net , \coefcal1_divide_inst1_u107_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_1|SUM_net , \coefcal1_divide_inst1_u107_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_3|SUM_net , \coefcal1_divide_inst1_u107_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_5|SUM_net , \coefcal1_divide_inst1_u107_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_7|SUM_net , \coefcal1_divide_inst1_u107_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u107_XORCI_9|SUM_net , \coefcal1_divide_inst1_u108_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_10|SUM_net , \coefcal1_divide_inst1_u108_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_12|SUM_net , \coefcal1_divide_inst1_u108_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_14|SUM_net , \coefcal1_divide_inst1_u108_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_1|SUM_net , \coefcal1_divide_inst1_u108_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_3|SUM_net , \coefcal1_divide_inst1_u108_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_5|SUM_net , \coefcal1_divide_inst1_u108_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_7|SUM_net , \coefcal1_divide_inst1_u108_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u108_XORCI_9|SUM_net , \coefcal1_divide_inst1_u109_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_10|SUM_net , \coefcal1_divide_inst1_u109_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_12|SUM_net , \coefcal1_divide_inst1_u109_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_14|SUM_net , \coefcal1_divide_inst1_u109_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_1|SUM_net , \coefcal1_divide_inst1_u109_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_3|SUM_net , \coefcal1_divide_inst1_u109_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_5|SUM_net , \coefcal1_divide_inst1_u109_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_7|SUM_net , \coefcal1_divide_inst1_u109_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u109_XORCI_9|SUM_net , \coefcal1_divide_inst1_u110_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_10|SUM_net , \coefcal1_divide_inst1_u110_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_12|SUM_net , \coefcal1_divide_inst1_u110_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_14|SUM_net , \coefcal1_divide_inst1_u110_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_1|SUM_net , \coefcal1_divide_inst1_u110_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_3|SUM_net , \coefcal1_divide_inst1_u110_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_5|SUM_net , \coefcal1_divide_inst1_u110_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_7|SUM_net , \coefcal1_divide_inst1_u110_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u110_XORCI_9|SUM_net , \coefcal1_divide_inst1_u111_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_10|SUM_net , \coefcal1_divide_inst1_u111_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_12|SUM_net , \coefcal1_divide_inst1_u111_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_14|SUM_net , \coefcal1_divide_inst1_u111_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_1|SUM_net , \coefcal1_divide_inst1_u111_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_3|SUM_net , \coefcal1_divide_inst1_u111_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_5|SUM_net , \coefcal1_divide_inst1_u111_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_7|SUM_net , \coefcal1_divide_inst1_u111_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u111_XORCI_9|SUM_net , \coefcal1_divide_inst1_u112_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_10|SUM_net , \coefcal1_divide_inst1_u112_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_12|SUM_net , \coefcal1_divide_inst1_u112_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_14|SUM_net , \coefcal1_divide_inst1_u112_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_1|SUM_net , \coefcal1_divide_inst1_u112_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_3|SUM_net , \coefcal1_divide_inst1_u112_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_5|SUM_net , \coefcal1_divide_inst1_u112_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_7|SUM_net , \coefcal1_divide_inst1_u112_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u112_XORCI_9|SUM_net , \coefcal1_divide_inst1_u113_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_10|SUM_net , \coefcal1_divide_inst1_u113_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_12|SUM_net , \coefcal1_divide_inst1_u113_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_14|SUM_net , \coefcal1_divide_inst1_u113_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_1|SUM_net , \coefcal1_divide_inst1_u113_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_3|SUM_net , \coefcal1_divide_inst1_u113_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_5|SUM_net , \coefcal1_divide_inst1_u113_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_7|SUM_net , \coefcal1_divide_inst1_u113_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u113_XORCI_9|SUM_net , \coefcal1_divide_inst1_u114_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_10|SUM_net , \coefcal1_divide_inst1_u114_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_12|SUM_net , \coefcal1_divide_inst1_u114_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_14|SUM_net , \coefcal1_divide_inst1_u114_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_1|SUM_net , \coefcal1_divide_inst1_u114_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_3|SUM_net , \coefcal1_divide_inst1_u114_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_5|SUM_net , \coefcal1_divide_inst1_u114_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_7|SUM_net , \coefcal1_divide_inst1_u114_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u114_XORCI_9|SUM_net , \coefcal1_divide_inst1_u115_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_10|SUM_net , \coefcal1_divide_inst1_u115_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_12|SUM_net , \coefcal1_divide_inst1_u115_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_14|SUM_net , \coefcal1_divide_inst1_u115_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_1|SUM_net , \coefcal1_divide_inst1_u115_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_3|SUM_net , \coefcal1_divide_inst1_u115_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_5|SUM_net , \coefcal1_divide_inst1_u115_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_7|SUM_net , \coefcal1_divide_inst1_u115_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u115_XORCI_9|SUM_net , \coefcal1_divide_inst1_u116_XORCI_0|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_10|SUM_net , \coefcal1_divide_inst1_u116_XORCI_11|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_12|SUM_net , \coefcal1_divide_inst1_u116_XORCI_13|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_14|SUM_net , \coefcal1_divide_inst1_u116_XORCI_15|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_1|SUM_net , \coefcal1_divide_inst1_u116_XORCI_2|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_3|SUM_net , \coefcal1_divide_inst1_u116_XORCI_4|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_5|SUM_net , \coefcal1_divide_inst1_u116_XORCI_6|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_7|SUM_net , \coefcal1_divide_inst1_u116_XORCI_8|SUM_net ,
       \coefcal1_divide_inst1_u116_XORCI_9|SUM_net , \coefcal1_divide_inst1_u118_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u120_XORCI_17|SUM_net , \coefcal1_divide_inst1_u122_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u124_XORCI_17|SUM_net , \coefcal1_divide_inst1_u126_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u128_XORCI_17|SUM_net , \coefcal1_divide_inst1_u130_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u132_XORCI_17|SUM_net , \coefcal1_divide_inst1_u134_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u136_XORCI_17|SUM_net , \coefcal1_divide_inst1_u138_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u140_XORCI_17|SUM_net , \coefcal1_divide_inst1_u142_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u144_XORCI_17|SUM_net , \coefcal1_divide_inst1_u146_XORCI_17|SUM_net ,
       \coefcal1_divide_inst1_u148_XORCI_17|SUM_net , \coefcal1_divide_inst1_u150_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_0|SUM_net , \coefcal1_divide_inst2_u102_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_11|SUM_net , \coefcal1_divide_inst2_u102_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_13|SUM_net , \coefcal1_divide_inst2_u102_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_15|SUM_net , \coefcal1_divide_inst2_u102_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_2|SUM_net , \coefcal1_divide_inst2_u102_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_4|SUM_net , \coefcal1_divide_inst2_u102_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_6|SUM_net , \coefcal1_divide_inst2_u102_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u102_XORCI_8|SUM_net , \coefcal1_divide_inst2_u102_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_0|SUM_net , \coefcal1_divide_inst2_u103_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_11|SUM_net , \coefcal1_divide_inst2_u103_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_13|SUM_net , \coefcal1_divide_inst2_u103_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_15|SUM_net , \coefcal1_divide_inst2_u103_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_2|SUM_net , \coefcal1_divide_inst2_u103_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_4|SUM_net , \coefcal1_divide_inst2_u103_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_6|SUM_net , \coefcal1_divide_inst2_u103_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u103_XORCI_8|SUM_net , \coefcal1_divide_inst2_u103_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_0|SUM_net , \coefcal1_divide_inst2_u104_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_11|SUM_net , \coefcal1_divide_inst2_u104_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_13|SUM_net , \coefcal1_divide_inst2_u104_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_15|SUM_net , \coefcal1_divide_inst2_u104_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_2|SUM_net , \coefcal1_divide_inst2_u104_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_4|SUM_net , \coefcal1_divide_inst2_u104_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_6|SUM_net , \coefcal1_divide_inst2_u104_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u104_XORCI_8|SUM_net , \coefcal1_divide_inst2_u104_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_0|SUM_net , \coefcal1_divide_inst2_u105_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_11|SUM_net , \coefcal1_divide_inst2_u105_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_13|SUM_net , \coefcal1_divide_inst2_u105_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_15|SUM_net , \coefcal1_divide_inst2_u105_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_2|SUM_net , \coefcal1_divide_inst2_u105_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_4|SUM_net , \coefcal1_divide_inst2_u105_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_6|SUM_net , \coefcal1_divide_inst2_u105_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u105_XORCI_8|SUM_net , \coefcal1_divide_inst2_u105_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_0|SUM_net , \coefcal1_divide_inst2_u106_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_11|SUM_net , \coefcal1_divide_inst2_u106_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_13|SUM_net , \coefcal1_divide_inst2_u106_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_15|SUM_net , \coefcal1_divide_inst2_u106_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_2|SUM_net , \coefcal1_divide_inst2_u106_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_4|SUM_net , \coefcal1_divide_inst2_u106_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_6|SUM_net , \coefcal1_divide_inst2_u106_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u106_XORCI_8|SUM_net , \coefcal1_divide_inst2_u106_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_0|SUM_net , \coefcal1_divide_inst2_u107_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_11|SUM_net , \coefcal1_divide_inst2_u107_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_13|SUM_net , \coefcal1_divide_inst2_u107_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_15|SUM_net , \coefcal1_divide_inst2_u107_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_2|SUM_net , \coefcal1_divide_inst2_u107_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_4|SUM_net , \coefcal1_divide_inst2_u107_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_6|SUM_net , \coefcal1_divide_inst2_u107_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u107_XORCI_8|SUM_net , \coefcal1_divide_inst2_u107_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_0|SUM_net , \coefcal1_divide_inst2_u108_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_11|SUM_net , \coefcal1_divide_inst2_u108_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_13|SUM_net , \coefcal1_divide_inst2_u108_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_15|SUM_net , \coefcal1_divide_inst2_u108_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_2|SUM_net , \coefcal1_divide_inst2_u108_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_4|SUM_net , \coefcal1_divide_inst2_u108_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_6|SUM_net , \coefcal1_divide_inst2_u108_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u108_XORCI_8|SUM_net , \coefcal1_divide_inst2_u108_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_0|SUM_net , \coefcal1_divide_inst2_u109_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_11|SUM_net , \coefcal1_divide_inst2_u109_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_13|SUM_net , \coefcal1_divide_inst2_u109_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_15|SUM_net , \coefcal1_divide_inst2_u109_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_2|SUM_net , \coefcal1_divide_inst2_u109_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_4|SUM_net , \coefcal1_divide_inst2_u109_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_6|SUM_net , \coefcal1_divide_inst2_u109_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u109_XORCI_8|SUM_net , \coefcal1_divide_inst2_u109_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_0|SUM_net , \coefcal1_divide_inst2_u110_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_11|SUM_net , \coefcal1_divide_inst2_u110_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_13|SUM_net , \coefcal1_divide_inst2_u110_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_15|SUM_net , \coefcal1_divide_inst2_u110_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_2|SUM_net , \coefcal1_divide_inst2_u110_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_4|SUM_net , \coefcal1_divide_inst2_u110_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_6|SUM_net , \coefcal1_divide_inst2_u110_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u110_XORCI_8|SUM_net , \coefcal1_divide_inst2_u110_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_0|SUM_net , \coefcal1_divide_inst2_u111_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_11|SUM_net , \coefcal1_divide_inst2_u111_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_13|SUM_net , \coefcal1_divide_inst2_u111_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_15|SUM_net , \coefcal1_divide_inst2_u111_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_2|SUM_net , \coefcal1_divide_inst2_u111_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_4|SUM_net , \coefcal1_divide_inst2_u111_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_6|SUM_net , \coefcal1_divide_inst2_u111_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u111_XORCI_8|SUM_net , \coefcal1_divide_inst2_u111_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_0|SUM_net , \coefcal1_divide_inst2_u112_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_11|SUM_net , \coefcal1_divide_inst2_u112_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_13|SUM_net , \coefcal1_divide_inst2_u112_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_15|SUM_net , \coefcal1_divide_inst2_u112_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_2|SUM_net , \coefcal1_divide_inst2_u112_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_4|SUM_net , \coefcal1_divide_inst2_u112_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_6|SUM_net , \coefcal1_divide_inst2_u112_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u112_XORCI_8|SUM_net , \coefcal1_divide_inst2_u112_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_0|SUM_net , \coefcal1_divide_inst2_u113_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_11|SUM_net , \coefcal1_divide_inst2_u113_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_13|SUM_net , \coefcal1_divide_inst2_u113_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_15|SUM_net , \coefcal1_divide_inst2_u113_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_2|SUM_net , \coefcal1_divide_inst2_u113_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_4|SUM_net , \coefcal1_divide_inst2_u113_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_6|SUM_net , \coefcal1_divide_inst2_u113_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u113_XORCI_8|SUM_net , \coefcal1_divide_inst2_u113_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_0|SUM_net , \coefcal1_divide_inst2_u114_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_11|SUM_net , \coefcal1_divide_inst2_u114_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_13|SUM_net , \coefcal1_divide_inst2_u114_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_15|SUM_net , \coefcal1_divide_inst2_u114_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_2|SUM_net , \coefcal1_divide_inst2_u114_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_4|SUM_net , \coefcal1_divide_inst2_u114_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_6|SUM_net , \coefcal1_divide_inst2_u114_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u114_XORCI_8|SUM_net , \coefcal1_divide_inst2_u114_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_0|SUM_net , \coefcal1_divide_inst2_u115_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_11|SUM_net , \coefcal1_divide_inst2_u115_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_13|SUM_net , \coefcal1_divide_inst2_u115_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_15|SUM_net , \coefcal1_divide_inst2_u115_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_2|SUM_net , \coefcal1_divide_inst2_u115_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_4|SUM_net , \coefcal1_divide_inst2_u115_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_6|SUM_net , \coefcal1_divide_inst2_u115_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u115_XORCI_8|SUM_net , \coefcal1_divide_inst2_u115_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_0|SUM_net , \coefcal1_divide_inst2_u116_XORCI_10|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_11|SUM_net , \coefcal1_divide_inst2_u116_XORCI_12|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_13|SUM_net , \coefcal1_divide_inst2_u116_XORCI_14|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_15|SUM_net , \coefcal1_divide_inst2_u116_XORCI_1|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_2|SUM_net , \coefcal1_divide_inst2_u116_XORCI_3|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_4|SUM_net , \coefcal1_divide_inst2_u116_XORCI_5|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_6|SUM_net , \coefcal1_divide_inst2_u116_XORCI_7|SUM_net ,
       \coefcal1_divide_inst2_u116_XORCI_8|SUM_net , \coefcal1_divide_inst2_u116_XORCI_9|SUM_net ,
       \coefcal1_divide_inst2_u118_XORCI_17|SUM_net , \coefcal1_divide_inst2_u120_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u122_XORCI_17|SUM_net , \coefcal1_divide_inst2_u124_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u126_XORCI_17|SUM_net , \coefcal1_divide_inst2_u128_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u130_XORCI_17|SUM_net , \coefcal1_divide_inst2_u132_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u134_XORCI_17|SUM_net , \coefcal1_divide_inst2_u136_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u138_XORCI_17|SUM_net , \coefcal1_divide_inst2_u140_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u142_XORCI_17|SUM_net , \coefcal1_divide_inst2_u144_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u146_XORCI_17|SUM_net , \coefcal1_divide_inst2_u148_XORCI_17|SUM_net ,
       \coefcal1_divide_inst2_u150_XORCI_17|SUM_net , \coefcal1_frameRate__reg[0]|Q_net ,
       \coefcal1_frameRate__reg[1]|Q_net , \coefcal1_frameRate__reg[2]|Q_net ,
       \coefcal1_frameRate__reg[3]|Q_net , \coefcal1_frameRate__reg[4]|Q_net ,
       \coefcal1_frameRate__reg[5]|Q_net , \coefcal1_frameRate__reg[6]|Q_net ,
       \coefcal1_frameRate__reg[7]|Q_net , \coefcal1_frameRate__reg[8]|Q_net ,
       \coefcal1_inEn__reg|Q_net , \coefcal1_u59_XORCI_0|SUM_net , \coefcal1_u59_XORCI_10|SUM_net ,
       \coefcal1_u59_XORCI_1|SUM_net , \coefcal1_u59_XORCI_2|SUM_net , \coefcal1_u59_XORCI_3|SUM_net ,
       \coefcal1_u59_XORCI_4|SUM_net , \coefcal1_u59_XORCI_5|SUM_net , \coefcal1_u59_XORCI_6|SUM_net ,
       \coefcal1_u59_XORCI_7|SUM_net , \coefcal1_u59_XORCI_8|SUM_net , \coefcal1_u59_XORCI_9|SUM_net ,
       \coefcal1_u60_XORCI_0|SUM_net , \coefcal1_u60_XORCI_10|SUM_net , \coefcal1_u60_XORCI_1|SUM_net ,
       \coefcal1_u60_XORCI_2|SUM_net , \coefcal1_u60_XORCI_3|SUM_net , \coefcal1_u60_XORCI_4|SUM_net ,
       \coefcal1_u60_XORCI_5|SUM_net , \coefcal1_u60_XORCI_6|SUM_net , \coefcal1_u60_XORCI_7|SUM_net ,
       \coefcal1_u60_XORCI_8|SUM_net , \coefcal1_u60_XORCI_9|SUM_net , \coefcal1_u61_XORCI_0|SUM_net ,
       \coefcal1_u61_XORCI_1|SUM_net , \coefcal1_u61_XORCI_2|SUM_net , \coefcal1_u61_XORCI_3|SUM_net ,
       \coefcal1_u61_XORCI_4|SUM_net , \coefcal1_u61_XORCI_5|SUM_net , \coefcal1_u61_XORCI_6|SUM_net ,
       \coefcal1_u61_XORCI_7|SUM_net , \coefcal1_u62_XORCI_0|SUM_net , \coefcal1_u62_XORCI_1|SUM_net ,
       \coefcal1_u62_XORCI_2|SUM_net , \coefcal1_u62_XORCI_3|SUM_net , \coefcal1_u62_XORCI_4|SUM_net ,
       \coefcal1_u62_XORCI_5|SUM_net , \coefcal1_u62_XORCI_6|SUM_net , \coefcal1_u62_XORCI_7|SUM_net ,
       \coefcal1_u64_XORCI_0|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , \coefcal1_u64_XORCI_11|SUM_net ,
       \coefcal1_u64_XORCI_12|SUM_net , \coefcal1_u64_XORCI_1|SUM_net , \coefcal1_u64_XORCI_2|SUM_net ,
       \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , \coefcal1_u64_XORCI_5|SUM_net ,
       \coefcal1_u64_XORCI_6|SUM_net , \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_8|SUM_net ,
       \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u7_XORCI_0|SUM_net , \coefcal1_u7_XORCI_10|SUM_net ,
       \coefcal1_u7_XORCI_1|SUM_net , \coefcal1_u7_XORCI_2|SUM_net , \coefcal1_u7_XORCI_3|SUM_net ,
       \coefcal1_u7_XORCI_4|SUM_net , \coefcal1_u7_XORCI_5|SUM_net , \coefcal1_u7_XORCI_6|SUM_net ,
       \coefcal1_u7_XORCI_7|SUM_net , \coefcal1_u7_XORCI_8|SUM_net , \coefcal1_u7_XORCI_9|SUM_net ,
       \coefcal1_u8_XORCI_33|SUM_net , \coefcal1_work__reg|Q_net , \coefcal1_working__reg[0]|Q_net ,
       \coefcal1_working__reg[10]|Q_net , \coefcal1_working__reg[11]|Q_net ,
       \coefcal1_working__reg[12]|Q_net , \coefcal1_working__reg[13]|Q_net ,
       \coefcal1_working__reg[14]|Q_net , \coefcal1_working__reg[15]|Q_net ,
       \coefcal1_working__reg[16]|Q_net , \coefcal1_working__reg[17]|Q_net ,
       \coefcal1_working__reg[18]|Q_net , \coefcal1_working__reg[19]|Q_net ,
       \coefcal1_working__reg[1]|Q_net , \coefcal1_working__reg[20]|Q_net , \coefcal1_working__reg[21]|Q_net ,
       \coefcal1_working__reg[22]|Q_net , \coefcal1_working__reg[23]|Q_net ,
       \coefcal1_working__reg[24]|Q_net , \coefcal1_working__reg[25]|Q_net ,
       \coefcal1_working__reg[26]|Q_net , \coefcal1_working__reg[27]|Q_net ,
       \coefcal1_working__reg[28]|Q_net , \coefcal1_working__reg[29]|Q_net ,
       \coefcal1_working__reg[2]|Q_net , \coefcal1_working__reg[30]|Q_net , \coefcal1_working__reg[31]|Q_net ,
       \coefcal1_working__reg[32]|Q_net , \coefcal1_working__reg[3]|Q_net , \coefcal1_working__reg[4]|Q_net ,
       \coefcal1_working__reg[5]|Q_net , \coefcal1_working__reg[6]|Q_net , \coefcal1_working__reg[7]|Q_net ,
       \coefcal1_working__reg[8]|Q_net , \coefcal1_working__reg[9]|Q_net , \coefcal1_xDividend__reg[0]|Q_net ,
       \coefcal1_xDividend__reg[10]|Q_net , \coefcal1_xDividend__reg[11]|Q_net ,
       \coefcal1_xDividend__reg[12]|Q_net , \coefcal1_xDividend__reg[13]|Q_net ,
       \coefcal1_xDividend__reg[14]|Q_net , \coefcal1_xDividend__reg[15]|Q_net ,
       \coefcal1_xDividend__reg[16]|Q_net , \coefcal1_xDividend__reg[1]|Q_net ,
       \coefcal1_xDividend__reg[2]|Q_net , \coefcal1_xDividend__reg[3]|Q_net ,
       \coefcal1_xDividend__reg[4]|Q_net , \coefcal1_xDividend__reg[5]|Q_net ,
       \coefcal1_xDividend__reg[6]|Q_net , \coefcal1_xDividend__reg[7]|Q_net ,
       \coefcal1_xDividend__reg[8]|Q_net , \coefcal1_xDividend__reg[9]|Q_net ,
       \coefcal1_xDivisor__reg[0]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net ,
       \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net ,
       \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net ,
       \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[16]|Q_net ,
       \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net ,
       \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net ,
       \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net ,
       \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net ,
       \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_yDividend__reg[0]|Q_net ,
       \coefcal1_yDividend__reg[10]|Q_net , \coefcal1_yDividend__reg[11]|Q_net ,
       \coefcal1_yDividend__reg[12]|Q_net , \coefcal1_yDividend__reg[13]|Q_net ,
       \coefcal1_yDividend__reg[14]|Q_net , \coefcal1_yDividend__reg[15]|Q_net ,
       \coefcal1_yDividend__reg[16]|Q_net , \coefcal1_yDividend__reg[1]|Q_net ,
       \coefcal1_yDividend__reg[2]|Q_net , \coefcal1_yDividend__reg[3]|Q_net ,
       \coefcal1_yDividend__reg[4]|Q_net , \coefcal1_yDividend__reg[5]|Q_net ,
       \coefcal1_yDividend__reg[6]|Q_net , \coefcal1_yDividend__reg[7]|Q_net ,
       \coefcal1_yDividend__reg[8]|Q_net , \coefcal1_yDividend__reg[9]|Q_net ,
       \coefcal1_yDivisor__reg[0]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net ,
       \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net ,
       \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net ,
       \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[16]|Q_net ,
       \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net ,
       \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net ,
       \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net ,
       \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net ,
       \coefcal1_yDivisor__reg[9]|Q_net , dOut_0__net, dOut_10__net, dOut_11__net,
       dOut_12__net, dOut_13__net, dOut_14__net, dOut_15__net, dOut_16__net,
       dOut_17__net, dOut_18__net, dOut_19__net, dOut_1__net, dOut_20__net, dOut_21__net,
       dOut_22__net, dOut_23__net, dOut_2__net, dOut_3__net, dOut_4__net, dOut_5__net,
       dOut_6__net, dOut_7__net, dOut_8__net, dOut_9__net, \fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_3A_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_3A_ab_reg__reg[0]|Q_net , \fifo1_ram_inst_3B_aa_reg__reg[0]|Q_net ,
       \fifo1_ram_inst_3B_ab_reg__reg[0]|Q_net , \inputctrl1_dataOut__reg[0]|Q_net ,
       \inputctrl1_dataOut__reg[10]|Q_net , \inputctrl1_dataOut__reg[11]|Q_net ,
       \inputctrl1_dataOut__reg[12]|Q_net , \inputctrl1_dataOut__reg[13]|Q_net ,
       \inputctrl1_dataOut__reg[14]|Q_net , \inputctrl1_dataOut__reg[15]|Q_net ,
       \inputctrl1_dataOut__reg[16]|Q_net , \inputctrl1_dataOut__reg[17]|Q_net ,
       \inputctrl1_dataOut__reg[18]|Q_net , \inputctrl1_dataOut__reg[19]|Q_net ,
       \inputctrl1_dataOut__reg[1]|Q_net , \inputctrl1_dataOut__reg[20]|Q_net ,
       \inputctrl1_dataOut__reg[21]|Q_net , \inputctrl1_dataOut__reg[22]|Q_net ,
       \inputctrl1_dataOut__reg[23]|Q_net , \inputctrl1_dataOut__reg[2]|Q_net ,
       \inputctrl1_dataOut__reg[3]|Q_net , \inputctrl1_dataOut__reg[4]|Q_net ,
       \inputctrl1_dataOut__reg[5]|Q_net , \inputctrl1_dataOut__reg[6]|Q_net ,
       \inputctrl1_dataOut__reg[7]|Q_net , \inputctrl1_dataOut__reg[8]|Q_net ,
       \inputctrl1_dataOut__reg[9]|Q_net , \inputctrl1_jmp__reg|Q_net , \inputctrl1_ramWrtAddr__reg[0]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[10]|Q_net , \inputctrl1_ramWrtAddr__reg[1]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[2]|Q_net , \inputctrl1_ramWrtAddr__reg[3]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[4]|Q_net , \inputctrl1_ramWrtAddr__reg[5]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[6]|Q_net , \inputctrl1_ramWrtAddr__reg[7]|Q_net ,
       \inputctrl1_ramWrtAddr__reg[8]|Q_net , \inputctrl1_ramWrtAddr__reg[9]|Q_net ,
       \inputctrl1_ramWrtEn__reg|Q_net , \inputctrl1_u108_XORCI_0|SUM_net , \inputctrl1_u108_XORCI_10|SUM_net ,
       \inputctrl1_u108_XORCI_11|SUM_net , \inputctrl1_u108_XORCI_12|SUM_net ,
       \inputctrl1_u108_XORCI_13|SUM_net , \inputctrl1_u108_XORCI_14|SUM_net ,
       \inputctrl1_u108_XORCI_15|SUM_net , \inputctrl1_u108_XORCI_16|SUM_net ,
       \inputctrl1_u108_XORCI_1|SUM_net , \inputctrl1_u108_XORCI_2|SUM_net ,
       \inputctrl1_u108_XORCI_3|SUM_net , \inputctrl1_u108_XORCI_4|SUM_net ,
       \inputctrl1_u108_XORCI_5|SUM_net , \inputctrl1_u108_XORCI_6|SUM_net ,
       \inputctrl1_u108_XORCI_7|SUM_net , \inputctrl1_u108_XORCI_8|SUM_net ,
       \inputctrl1_u108_XORCI_9|SUM_net , \inputctrl1_u109_XORCI_0|SUM_net ,
       \inputctrl1_u109_XORCI_10|SUM_net , \inputctrl1_u109_XORCI_11|SUM_net ,
       \inputctrl1_u109_XORCI_12|SUM_net , \inputctrl1_u109_XORCI_13|SUM_net ,
       \inputctrl1_u109_XORCI_14|SUM_net , \inputctrl1_u109_XORCI_15|SUM_net ,
       \inputctrl1_u109_XORCI_16|SUM_net , \inputctrl1_u109_XORCI_1|SUM_net ,
       \inputctrl1_u109_XORCI_2|SUM_net , \inputctrl1_u109_XORCI_3|SUM_net ,
       \inputctrl1_u109_XORCI_4|SUM_net , \inputctrl1_u109_XORCI_5|SUM_net ,
       \inputctrl1_u109_XORCI_6|SUM_net , \inputctrl1_u109_XORCI_7|SUM_net ,
       \inputctrl1_u109_XORCI_8|SUM_net , \inputctrl1_u109_XORCI_9|SUM_net ,
       \inputctrl1_u110_XORCI_0|SUM_net , \inputctrl1_u110_XORCI_10|SUM_net ,
       \inputctrl1_u110_XORCI_1|SUM_net , \inputctrl1_u110_XORCI_2|SUM_net ,
       \inputctrl1_u110_XORCI_3|SUM_net , \inputctrl1_u110_XORCI_4|SUM_net ,
       \inputctrl1_u110_XORCI_5|SUM_net , \inputctrl1_u110_XORCI_6|SUM_net ,
       \inputctrl1_u110_XORCI_7|SUM_net , \inputctrl1_u110_XORCI_8|SUM_net ,
       \inputctrl1_u110_XORCI_9|SUM_net , \inputctrl1_u111_XORCI_0|SUM_net ,
       \inputctrl1_u111_XORCI_10|SUM_net , \inputctrl1_u111_XORCI_1|SUM_net ,
       \inputctrl1_u111_XORCI_2|SUM_net , \inputctrl1_u111_XORCI_3|SUM_net ,
       \inputctrl1_u111_XORCI_4|SUM_net , \inputctrl1_u111_XORCI_5|SUM_net ,
       \inputctrl1_u111_XORCI_6|SUM_net , \inputctrl1_u111_XORCI_7|SUM_net ,
       \inputctrl1_u111_XORCI_8|SUM_net , \inputctrl1_u111_XORCI_9|SUM_net ,
       \inputctrl1_u112_XORCI_0|SUM_net , \inputctrl1_u112_XORCI_10|SUM_net ,
       \inputctrl1_u112_XORCI_1|SUM_net , \inputctrl1_u112_XORCI_2|SUM_net ,
       \inputctrl1_u112_XORCI_3|SUM_net , \inputctrl1_u112_XORCI_4|SUM_net ,
       \inputctrl1_u112_XORCI_5|SUM_net , \inputctrl1_u112_XORCI_6|SUM_net ,
       \inputctrl1_u112_XORCI_7|SUM_net , \inputctrl1_u112_XORCI_8|SUM_net ,
       \inputctrl1_u112_XORCI_9|SUM_net , \inputctrl1_u37_XORCI_11|SUM_net ,
       \inputctrl1_u39_XORCI_11|SUM_net , \inputctrl1_u41_XORCI_11|SUM_net ,
       \inputctrl1_u43_XORCI_11|SUM_net , \inputctrl1_xAddress__reg[0]|Q_net ,
       \inputctrl1_xAddress__reg[10]|Q_net , \inputctrl1_xAddress__reg[1]|Q_net ,
       \inputctrl1_xAddress__reg[2]|Q_net , \inputctrl1_xAddress__reg[3]|Q_net ,
       \inputctrl1_xAddress__reg[4]|Q_net , \inputctrl1_xAddress__reg[5]|Q_net ,
       \inputctrl1_xAddress__reg[6]|Q_net , \inputctrl1_xAddress__reg[7]|Q_net ,
       \inputctrl1_xAddress__reg[8]|Q_net , \inputctrl1_xAddress__reg[9]|Q_net ,
       \inputctrl1_xCal__reg[0]|Q_net , \inputctrl1_xCal__reg[10]|Q_net , \inputctrl1_xCal__reg[11]|Q_net ,
       \inputctrl1_xCal__reg[12]|Q_net , \inputctrl1_xCal__reg[13]|Q_net , \inputctrl1_xCal__reg[14]|Q_net ,
       \inputctrl1_xCal__reg[15]|Q_net , \inputctrl1_xCal__reg[16]|Q_net , \inputctrl1_xCal__reg[1]|Q_net ,
       \inputctrl1_xCal__reg[2]|Q_net , \inputctrl1_xCal__reg[3]|Q_net , \inputctrl1_xCal__reg[4]|Q_net ,
       \inputctrl1_xCal__reg[5]|Q_net , \inputctrl1_xCal__reg[6]|Q_net , \inputctrl1_xCal__reg[7]|Q_net ,
       \inputctrl1_xCal__reg[8]|Q_net , \inputctrl1_xCal__reg[9]|Q_net , \inputctrl1_xPreEn__reg|Q_net ,
       \inputctrl1_yAddress__reg[0]|Q_net , \inputctrl1_yAddress__reg[10]|Q_net ,
       \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net ,
       \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net ,
       \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net ,
       \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net ,
       \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yCal__reg[0]|Q_net ,
       \inputctrl1_yCal__reg[10]|Q_net , \inputctrl1_yCal__reg[11]|Q_net , \inputctrl1_yCal__reg[12]|Q_net ,
       \inputctrl1_yCal__reg[13]|Q_net , \inputctrl1_yCal__reg[14]|Q_net , \inputctrl1_yCal__reg[15]|Q_net ,
       \inputctrl1_yCal__reg[16]|Q_net , \inputctrl1_yCal__reg[1]|Q_net , \inputctrl1_yCal__reg[2]|Q_net ,
       \inputctrl1_yCal__reg[3]|Q_net , \inputctrl1_yCal__reg[4]|Q_net , \inputctrl1_yCal__reg[5]|Q_net ,
       \inputctrl1_yCal__reg[6]|Q_net , \inputctrl1_yCal__reg[7]|Q_net , \inputctrl1_yCal__reg[8]|Q_net ,
       \inputctrl1_yCal__reg[9]|Q_net , \inputctrl1_yPreEn__reg|Q_net , \u2_XORCI_0|SUM_net ,
       \u2_XORCI_10|SUM_net , \u2_XORCI_11|SUM_net , \u2_XORCI_1|SUM_net , \u2_XORCI_2|SUM_net ,
       \u2_XORCI_3|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_5|SUM_net , \u2_XORCI_6|SUM_net ,
       \u2_XORCI_7|SUM_net , \u2_XORCI_8|SUM_net , \u2_XORCI_9|SUM_net , \u3_XORCI_0|SUM_net ,
       \u3_XORCI_10|SUM_net , \u3_XORCI_1|SUM_net , \u3_XORCI_2|SUM_net , \u3_XORCI_3|SUM_net ,
       \u3_XORCI_4|SUM_net , \u3_XORCI_5|SUM_net , \u3_XORCI_6|SUM_net , \u3_XORCI_7|SUM_net ,
       \u3_XORCI_8|SUM_net , \u3_XORCI_9|SUM_net ;

    assign HS = HS_2079_net;
    assign a_acc_en_cal1_u138_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u139_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u140_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u141_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u142_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u143_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u144_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u145_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u146_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u147_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u148_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_cal1_u149_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_coefcal1_u63_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign a_acc_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign \a_dinx[0]_cal1_u137_mac  = \cal1_uPreF__reg[0]|Q_net ;
    assign \a_dinx[0]_coefcal1_u63_mac  = outYRes[0];
    assign \a_dinx[0]_coefcal1_u64_mac  = \a_mac_out[0]_coefcal1_u63_mac ;
    assign \a_dinx[0]_coefcal1_u64_mac_0_  = \a_mac_out[18]_coefcal1_u63_mac ;
    assign \a_dinx[10]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_coefcal1_u63_mac  = outYRes[10];
    assign \a_dinx[10]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[10]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_coefcal1_u63_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[11]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_coefcal1_u63_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[12]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_coefcal1_u63_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[13]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[1]_cal1_u137_mac  = \cal1_uPreF__reg[1]|Q_net ;
    assign \a_dinx[1]_coefcal1_u63_mac  = outYRes[1];
    assign \a_dinx[1]_coefcal1_u64_mac  = \a_mac_out[1]_coefcal1_u63_mac ;
    assign \a_dinx[1]_coefcal1_u64_mac_0_  = \a_mac_out[19]_coefcal1_u63_mac ;
    assign \a_dinx[2]_cal1_u137_mac  = \cal1_uPreF__reg[2]|Q_net ;
    assign \a_dinx[2]_coefcal1_u63_mac  = outYRes[2];
    assign \a_dinx[2]_coefcal1_u64_mac  = \a_mac_out[2]_coefcal1_u63_mac ;
    assign \a_dinx[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[3]_cal1_u137_mac  = \cal1_uPreF__reg[3]|Q_net ;
    assign \a_dinx[3]_coefcal1_u63_mac  = outYRes[3];
    assign \a_dinx[3]_coefcal1_u64_mac  = \a_mac_out[3]_coefcal1_u63_mac ;
    assign \a_dinx[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[4]_cal1_u137_mac  = \cal1_uPreF__reg[4]|Q_net ;
    assign \a_dinx[4]_coefcal1_u63_mac  = outYRes[4];
    assign \a_dinx[4]_coefcal1_u64_mac  = \a_mac_out[4]_coefcal1_u63_mac ;
    assign \a_dinx[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[5]_cal1_u137_mac  = \cal1_uPreF__reg[5]|Q_net ;
    assign \a_dinx[5]_coefcal1_u63_mac  = outYRes[5];
    assign \a_dinx[5]_coefcal1_u64_mac  = \a_mac_out[5]_coefcal1_u63_mac ;
    assign \a_dinx[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[6]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[6]_coefcal1_u63_mac  = outYRes[6];
    assign \a_dinx[6]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[7]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[7]_coefcal1_u63_mac  = outYRes[7];
    assign \a_dinx[7]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_coefcal1_u63_mac  = outYRes[8];
    assign \a_dinx[8]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_coefcal1_u63_mac  = outYRes[9];
    assign \a_dinx[9]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_dinx[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u138_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u139_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u140_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u141_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u142_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u143_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u144_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u145_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u146_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u147_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u148_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_cal1_u149_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinxy_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign \a_diny[0]_cal1_u137_mac  = \cal1_v__reg[0]|Q_net ;
    assign \a_diny[0]_cal1_u138_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_diny[0]_cal1_u141_mac  = \a_mac_out[6]_cal1_u137_mac ;
    assign \a_diny[0]_cal1_u142_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_diny[0]_cal1_u143_mac  = \a_diny[0]_cal1_u139_mac ;
    assign \a_diny[0]_cal1_u144_mac  = \a_diny[0]_cal1_u140_mac ;
    assign \a_diny[0]_cal1_u145_mac  = \a_mac_out[6]_cal1_u137_mac ;
    assign \a_diny[0]_cal1_u146_mac  = \cal1_u133_XORCI_0|SUM_net ;
    assign \a_diny[0]_cal1_u147_mac  = \a_diny[0]_cal1_u139_mac ;
    assign \a_diny[0]_cal1_u148_mac  = \a_diny[0]_cal1_u140_mac ;
    assign \a_diny[0]_cal1_u149_mac  = \a_mac_out[6]_cal1_u137_mac ;
    assign \a_diny[0]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[0]|Q_net ;
    assign \a_diny[0]_coefcal1_u64_mac  = outXRes[0];
    assign \a_diny[0]_coefcal1_u64_mac_0_  = outXRes[0];
    assign \a_diny[1]_cal1_u137_mac  = \cal1_v__reg[1]|Q_net ;
    assign \a_diny[1]_cal1_u138_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_diny[1]_cal1_u141_mac  = \a_mac_out[7]_cal1_u137_mac ;
    assign \a_diny[1]_cal1_u142_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_diny[1]_cal1_u143_mac  = \a_diny[1]_cal1_u139_mac ;
    assign \a_diny[1]_cal1_u144_mac  = \a_diny[1]_cal1_u140_mac ;
    assign \a_diny[1]_cal1_u145_mac  = \a_mac_out[7]_cal1_u137_mac ;
    assign \a_diny[1]_cal1_u146_mac  = \cal1_u133_XORCI_1|SUM_net ;
    assign \a_diny[1]_cal1_u147_mac  = \a_diny[1]_cal1_u139_mac ;
    assign \a_diny[1]_cal1_u148_mac  = \a_diny[1]_cal1_u140_mac ;
    assign \a_diny[1]_cal1_u149_mac  = \a_mac_out[7]_cal1_u137_mac ;
    assign \a_diny[1]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[1]|Q_net ;
    assign \a_diny[1]_coefcal1_u64_mac  = outXRes[1];
    assign \a_diny[1]_coefcal1_u64_mac_0_  = outXRes[1];
    assign \a_diny[2]_cal1_u137_mac  = \cal1_v__reg[2]|Q_net ;
    assign \a_diny[2]_cal1_u138_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_diny[2]_cal1_u141_mac  = \a_mac_out[8]_cal1_u137_mac ;
    assign \a_diny[2]_cal1_u142_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_diny[2]_cal1_u143_mac  = \a_diny[2]_cal1_u139_mac ;
    assign \a_diny[2]_cal1_u144_mac  = \a_diny[2]_cal1_u140_mac ;
    assign \a_diny[2]_cal1_u145_mac  = \a_mac_out[8]_cal1_u137_mac ;
    assign \a_diny[2]_cal1_u146_mac  = \cal1_u133_XORCI_2|SUM_net ;
    assign \a_diny[2]_cal1_u147_mac  = \a_diny[2]_cal1_u139_mac ;
    assign \a_diny[2]_cal1_u148_mac  = \a_diny[2]_cal1_u140_mac ;
    assign \a_diny[2]_cal1_u149_mac  = \a_mac_out[8]_cal1_u137_mac ;
    assign \a_diny[2]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[2]|Q_net ;
    assign \a_diny[2]_coefcal1_u64_mac  = outXRes[2];
    assign \a_diny[2]_coefcal1_u64_mac_0_  = outXRes[2];
    assign \a_diny[3]_cal1_u137_mac  = \cal1_v__reg[3]|Q_net ;
    assign \a_diny[3]_cal1_u138_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_diny[3]_cal1_u141_mac  = \a_mac_out[9]_cal1_u137_mac ;
    assign \a_diny[3]_cal1_u142_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_diny[3]_cal1_u143_mac  = \a_diny[3]_cal1_u139_mac ;
    assign \a_diny[3]_cal1_u144_mac  = \a_diny[3]_cal1_u140_mac ;
    assign \a_diny[3]_cal1_u145_mac  = \a_mac_out[9]_cal1_u137_mac ;
    assign \a_diny[3]_cal1_u146_mac  = \cal1_u133_XORCI_3|SUM_net ;
    assign \a_diny[3]_cal1_u147_mac  = \a_diny[3]_cal1_u139_mac ;
    assign \a_diny[3]_cal1_u148_mac  = \a_diny[3]_cal1_u140_mac ;
    assign \a_diny[3]_cal1_u149_mac  = \a_mac_out[9]_cal1_u137_mac ;
    assign \a_diny[3]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[3]|Q_net ;
    assign \a_diny[3]_coefcal1_u64_mac  = outXRes[3];
    assign \a_diny[3]_coefcal1_u64_mac_0_  = outXRes[3];
    assign \a_diny[4]_cal1_u137_mac  = \cal1_v__reg[4]|Q_net ;
    assign \a_diny[4]_cal1_u138_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_diny[4]_cal1_u141_mac  = \a_mac_out[10]_cal1_u137_mac ;
    assign \a_diny[4]_cal1_u142_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_diny[4]_cal1_u143_mac  = \a_diny[4]_cal1_u139_mac ;
    assign \a_diny[4]_cal1_u144_mac  = \a_diny[4]_cal1_u140_mac ;
    assign \a_diny[4]_cal1_u145_mac  = \a_mac_out[10]_cal1_u137_mac ;
    assign \a_diny[4]_cal1_u146_mac  = \cal1_u133_XORCI_4|SUM_net ;
    assign \a_diny[4]_cal1_u147_mac  = \a_diny[4]_cal1_u139_mac ;
    assign \a_diny[4]_cal1_u148_mac  = \a_diny[4]_cal1_u140_mac ;
    assign \a_diny[4]_cal1_u149_mac  = \a_mac_out[10]_cal1_u137_mac ;
    assign \a_diny[4]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[4]|Q_net ;
    assign \a_diny[4]_coefcal1_u64_mac  = outXRes[4];
    assign \a_diny[4]_coefcal1_u64_mac_0_  = outXRes[4];
    assign \a_diny[5]_cal1_u137_mac  = \cal1_v__reg[5]|Q_net ;
    assign \a_diny[5]_cal1_u138_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_diny[5]_cal1_u141_mac  = \a_mac_out[11]_cal1_u137_mac ;
    assign \a_diny[5]_cal1_u142_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_diny[5]_cal1_u143_mac  = \a_diny[5]_cal1_u139_mac ;
    assign \a_diny[5]_cal1_u144_mac  = \a_diny[5]_cal1_u140_mac ;
    assign \a_diny[5]_cal1_u145_mac  = \a_mac_out[11]_cal1_u137_mac ;
    assign \a_diny[5]_cal1_u146_mac  = \cal1_u133_XORCI_5|SUM_net ;
    assign \a_diny[5]_cal1_u147_mac  = \a_diny[5]_cal1_u139_mac ;
    assign \a_diny[5]_cal1_u148_mac  = \a_diny[5]_cal1_u140_mac ;
    assign \a_diny[5]_cal1_u149_mac  = \a_mac_out[11]_cal1_u137_mac ;
    assign \a_diny[5]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[5]|Q_net ;
    assign \a_diny[5]_coefcal1_u64_mac  = outXRes[5];
    assign \a_diny[5]_coefcal1_u64_mac_0_  = outXRes[5];
    assign \a_diny[6]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u138_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_diny[6]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u142_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_diny[6]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u146_mac  = \cal1_u133_XORCI_6|SUM_net ;
    assign \a_diny[6]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[6]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[6]|Q_net ;
    assign \a_diny[6]_coefcal1_u64_mac  = outXRes[6];
    assign \a_diny[6]_coefcal1_u64_mac_0_  = outXRes[6];
    assign \a_diny[7]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[7]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[7]|Q_net ;
    assign \a_diny[7]_coefcal1_u64_mac  = outXRes[7];
    assign \a_diny[7]_coefcal1_u64_mac_0_  = outXRes[7];
    assign \a_diny[8]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[8]_coefcal1_u63_mac  = \coefcal1_frameRate__reg[8]|Q_net ;
    assign \a_diny[8]_coefcal1_u64_mac  = outXRes[8];
    assign \a_diny[8]_coefcal1_u64_mac_0_  = outXRes[8];
    assign \a_diny[9]_cal1_u137_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u138_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u139_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u140_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u141_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u142_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u143_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u144_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u145_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u146_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u147_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u148_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_cal1_u149_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_coefcal1_u63_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \a_diny[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign a_dinz_cen_cal1_u137_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u138_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u139_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u140_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u141_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u142_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u143_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u144_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u145_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u146_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u147_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u148_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_cal1_u149_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign a_dinz_en_cal1_u137_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u138_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u139_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u140_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u141_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u142_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u143_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u144_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u145_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u146_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u147_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u148_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_cal1_u149_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_coefcal1_u63_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign a_dinz_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign a_in_sr_cal1_u137_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u138_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u139_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u140_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u141_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u142_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u143_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u144_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u145_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u146_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u147_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u148_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_cal1_u149_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_coefcal1_u63_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_in_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u137_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u138_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u139_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u140_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u141_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u142_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u143_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u144_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u145_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u146_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u147_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u148_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_cal1_u149_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_coefcal1_u63_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_mac_out_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u137_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u138_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u139_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u140_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u141_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u142_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u143_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u144_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u145_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u146_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u147_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u148_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_cal1_u149_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_coefcal1_u63_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign a_out_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign a_sload_cal1_u137_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u138_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u139_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u140_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u141_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u142_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u143_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u144_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u145_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u146_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u147_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u148_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_cal1_u149_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_coefcal1_u63_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign a_sload_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign b_acc_en_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign b_acc_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign \b_dinx[0]_coefcal1_u64_mac  = \a_mac_out[6]_coefcal1_u63_mac ;
    assign \b_dinx[0]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[10]_coefcal1_u64_mac  = \a_mac_out[16]_coefcal1_u63_mac ;
    assign \b_dinx[10]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[11]_coefcal1_u64_mac  = \a_mac_out[17]_coefcal1_u63_mac ;
    assign \b_dinx[11]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[12]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[12]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[13]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[13]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[1]_coefcal1_u64_mac  = \a_mac_out[7]_coefcal1_u63_mac ;
    assign \b_dinx[1]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[2]_coefcal1_u64_mac  = \a_mac_out[8]_coefcal1_u63_mac ;
    assign \b_dinx[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[3]_coefcal1_u64_mac  = \a_mac_out[9]_coefcal1_u63_mac ;
    assign \b_dinx[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[4]_coefcal1_u64_mac  = \a_mac_out[10]_coefcal1_u63_mac ;
    assign \b_dinx[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[5]_coefcal1_u64_mac  = \a_mac_out[11]_coefcal1_u63_mac ;
    assign \b_dinx[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[6]_coefcal1_u64_mac  = \a_mac_out[12]_coefcal1_u63_mac ;
    assign \b_dinx[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[7]_coefcal1_u64_mac  = \a_mac_out[13]_coefcal1_u63_mac ;
    assign \b_dinx[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[8]_coefcal1_u64_mac  = \a_mac_out[14]_coefcal1_u63_mac ;
    assign \b_dinx[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_dinx[9]_coefcal1_u64_mac  = \a_mac_out[15]_coefcal1_u63_mac ;
    assign \b_dinx[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign b_dinxy_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign b_dinxy_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign \b_diny[0]_coefcal1_u64_mac  = outXRes[9];
    assign \b_diny[0]_coefcal1_u64_mac_0_  = outXRes[9];
    assign \b_diny[1]_coefcal1_u64_mac  = outXRes[10];
    assign \b_diny[1]_coefcal1_u64_mac_0_  = outXRes[10];
    assign \b_diny[2]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[2]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[3]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[3]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[4]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[4]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[5]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[5]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[6]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[6]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[7]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[7]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[8]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[8]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign \b_diny[9]_coefcal1_u64_mac  = a_acc_en_cal1_u137_mac;
    assign \b_diny[9]_coefcal1_u64_mac_0_  = a_acc_en_cal1_u137_mac;
    assign b_dinz_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign b_dinz_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign b_dinz_en_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign b_dinz_en_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign b_in_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign b_in_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign b_mac_out_cen_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign b_mac_out_cen_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign b_out_sr_coefcal1_u64_mac = a_dinxy_cen_cal1_u137_mac;
    assign b_out_sr_coefcal1_u64_mac_0_ = a_dinxy_cen_cal1_u137_mac;
    assign b_sload_coefcal1_u64_mac = a_acc_en_cal1_u137_mac;
    assign b_sload_coefcal1_u64_mac_0_ = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[10]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[11]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[2]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[3]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[4]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[5]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[6]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[7]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[8]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_0B_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_1B_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_2A_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_2B_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3A_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_0  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_aa[9]_fifo1_ram_inst_3B_u_emb18k_1  = \c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[10]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_8|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[11]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_9|SUM_net ;
    assign \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[2]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_0|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[3]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_1|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[4]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_2|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[5]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_3|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[6]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_4|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[7]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_5|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[8]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_6|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_7|SUM_net ;
    assign \c1r1_ab[9]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_7|SUM_net ;
    assign c1r1_clka_fifo1_ram_inst_0A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_0B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_0B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_1A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_1B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_1B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_2B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clka_fifo1_ram_inst_3B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_0A_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_0B_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1A_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_1B_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2A_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_2B_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3A_u_emb18k_1 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_0 = clkb;
    assign c1r1_clkb_fifo1_ram_inst_3B_u_emb18k_1 = clkb;
    assign \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[0]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[10]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[11]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[12]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[13]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[14]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[15]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[1]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[2]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[3]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[4]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[5]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r1_da[6]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r1_da[7]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r1_da[8]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r1_da[9]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r1_db[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstna_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r1_rstnb_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_clka_fifo1_ram_inst_0A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_0A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_0B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_0B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_1B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_2B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clka_fifo1_ram_inst_3B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_0A_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_0B_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1A_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_1B_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2A_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_2B_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3A_u_emb18k_1 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_0 = clkb;
    assign c1r2_clkb_fifo1_ram_inst_3B_u_emb18k_1 = clkb;
    assign \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r2_da[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r2_da[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r2_da[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r2_da[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r2_db[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstna_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r2_rstnb_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_clka_fifo1_ram_inst_0A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_0A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_0B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_0B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_1B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_2B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clka_fifo1_ram_inst_3B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_0A_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_0B_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1A_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_1B_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2A_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_2B_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3A_u_emb18k_1 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_0 = clkb;
    assign c1r3_clkb_fifo1_ram_inst_3B_u_emb18k_1 = clkb;
    assign \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[0]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[10]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[11]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[12]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[13]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[14]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[15]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[1]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[2]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[3]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[4]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[5]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[18]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[20]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[6]|Q_net ;
    assign \c1r3_da[6]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[8]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[21]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[23]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[9]|Q_net ;
    assign \c1r3_da[7]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[11]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[12]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[14]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[0]|Q_net ;
    assign \c1r3_da[8]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[2]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_0B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_1B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_2B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[15]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3A_u_emb18k_1  = \inputctrl1_dataOut__reg[17]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[3]|Q_net ;
    assign \c1r3_da[9]_fifo1_ram_inst_3B_u_emb18k_1  = \inputctrl1_dataOut__reg[5]|Q_net ;
    assign \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r3_db[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstna_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r3_rstnb_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_clka_fifo1_ram_inst_0A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_0A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_0B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_0B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_1B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_2B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3A_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3A_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3B_u_emb18k_0 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clka_fifo1_ram_inst_3B_u_emb18k_1 = c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0;
    assign c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_0A_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_0B_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1A_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_1B_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2A_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_2B_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3A_u_emb18k_1 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_0 = clkb;
    assign c1r4_clkb_fifo1_ram_inst_3B_u_emb18k_1 = clkb;
    assign \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[19]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[7]|Q_net ;
    assign \c1r4_da[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[22]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[10]|Q_net ;
    assign \c1r4_da[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[13]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[1]|Q_net ;
    assign \c1r4_da[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_0  = \inputctrl1_dataOut__reg[16]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_0  = \inputctrl1_dataOut__reg[4]|Q_net ;
    assign \c1r4_da[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[0]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[10]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[11]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[12]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[13]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[14]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[15]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[16]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[17]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[2]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[3]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[4]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[5]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[6]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[7]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[8]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \c1r4_db[9]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstna_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign c1r4_rstnb_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign cea_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_0A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_0A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_0B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_0B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_1A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_1A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_1B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_1B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_2A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_2A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_2B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_2B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_3A_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_3A_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_3B_u_emb18k_0 = a_dinxy_cen_cal1_u137_mac;
    assign ceb_fifo1_ram_inst_3B_u_emb18k_1 = a_dinxy_cen_cal1_u137_mac;
    assign dOut[0] = dOut_0__net;
    assign dOut[1] = dOut_1__net;
    assign dOut[2] = dOut_2__net;
    assign dOut[3] = dOut_3__net;
    assign dOut[4] = dOut_4__net;
    assign dOut[5] = dOut_5__net;
    assign dOut[6] = dOut_6__net;
    assign dOut[7] = dOut_7__net;
    assign dOut[8] = dOut_8__net;
    assign dOut[9] = dOut_9__net;
    assign dOut[10] = dOut_10__net;
    assign dOut[11] = dOut_11__net;
    assign dOut[12] = dOut_12__net;
    assign dOut[13] = dOut_13__net;
    assign dOut[14] = dOut_14__net;
    assign dOut[15] = dOut_15__net;
    assign dOut[16] = dOut_16__net;
    assign dOut[17] = dOut_17__net;
    assign dOut[18] = dOut_18__net;
    assign dOut[19] = dOut_19__net;
    assign dOut[20] = dOut_20__net;
    assign dOut[21] = dOut_21__net;
    assign dOut[22] = dOut_22__net;
    assign dOut[23] = dOut_23__net;
    assign \haa[0]_fifo1_ram_inst_0A_u_emb18k_1  = \haa[0]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_0B_u_emb18k_0  = \haa[0]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_0B_u_emb18k_1  = \haa[0]_fifo1_ram_inst_0A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_1A_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_1B_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_1B_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_2A_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_2A_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_2B_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_2B_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3A_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3A_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3B_u_emb18k_0  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[0]_fifo1_ram_inst_3B_u_emb18k_1  = \haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ;
    assign \haa[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \haa[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[0]_fifo1_ram_inst_0A_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_0A_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_0B_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_0B_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1A_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1A_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1B_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_1B_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2A_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2A_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2B_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_2B_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3A_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3A_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3B_u_emb18k_0  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[0]_fifo1_ram_inst_3B_u_emb18k_1  = \cal1_u129_XORCI_10|SUM_net ;
    assign \hab[1]_fifo1_ram_inst_0A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_0A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_0B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_0B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_1A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_1A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_1B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_1B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_2A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_2A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_2B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_2B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_3A_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_3A_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_3B_u_emb18k_0  = a_acc_en_cal1_u137_mac;
    assign \hab[1]_fifo1_ram_inst_3B_u_emb18k_1  = a_acc_en_cal1_u137_mac;
    assign u8205_O_1_ = u8205_O;
    assign u8205_O_2_ = u8205_O;
    assign u8224_O_4_ = u8224_O;
    assign wea_fifo1_ram_inst_0A_u_emb18k_1 = wea_fifo1_ram_inst_0A_u_emb18k_0;
    assign wea_fifo1_ram_inst_0B_u_emb18k_0 = wea_fifo1_ram_inst_0A_u_emb18k_0;
    assign wea_fifo1_ram_inst_0B_u_emb18k_1 = wea_fifo1_ram_inst_0A_u_emb18k_0;
    assign wea_fifo1_ram_inst_1A_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_1B_u_emb18k_0 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_1B_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_2A_u_emb18k_0 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_2A_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_2B_u_emb18k_0 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_2B_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_3A_u_emb18k_0 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_3A_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_3B_u_emb18k_0 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign wea_fifo1_ram_inst_3B_u_emb18k_1 = wea_fifo1_ram_inst_1A_u_emb18k_0;
    assign web_fifo1_ram_inst_0A_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_0A_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_0B_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_0B_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_1A_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_1A_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_1B_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_1B_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_2A_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_2A_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_2B_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_2B_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_3A_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_3A_u_emb18k_1 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_3B_u_emb18k_0 = a_acc_en_cal1_u137_mac;
    assign web_fifo1_ram_inst_3B_u_emb18k_1 = a_acc_en_cal1_u137_mac;

    CS_LUT4_PRIM ii0880 ( .DX(VS), .F0(\cal1_VSNormal__reg|Q_net ), .F1(\cal1_enforceJmp__reg|Q_net ), .F2(dummy_abc_1_), .F3(dummy_abc_2_) );
      defparam ii0880.CONFIG_DATA = 16'hEEEE;
      defparam ii0880.PLACE_LOCATION = "NONE";
      defparam ii0880.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0881 ( .DX(a_acc_en_cal1_u137_mac), .F0(dummy_abc_3_), .F1(dummy_abc_4_), .F2(dummy_abc_5_), .F3(dummy_abc_6_) );
      defparam ii0881.CONFIG_DATA = 16'h0000;
      defparam ii0881.PLACE_LOCATION = "NONE";
      defparam ii0881.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0882 ( .DX(nn0882), .F0(rst), .F1(u5502_IN), .F2(dummy_abc_7_), .F3(dummy_abc_8_) );
      defparam ii0882.CONFIG_DATA = 16'h2222;
      defparam ii0882.PLACE_LOCATION = "NONE";
      defparam ii0882.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0883 ( .DX(\a_dinx[0]_cal1_u138_mac ), .F0(\c1r2_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0883.CONFIG_DATA = 16'hCA00;
      defparam ii0883.PLACE_LOCATION = "NONE";
      defparam ii0883.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0884 ( .DX(\a_dinx[0]_cal1_u139_mac ), .F0(\c1r2_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0884.CONFIG_DATA = 16'hCA00;
      defparam ii0884.PLACE_LOCATION = "NONE";
      defparam ii0884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0885 ( .DX(a_dinxy_cen_cal1_u137_mac), .F0(dummy_abc_9_), .F1(dummy_abc_10_), .F2(dummy_abc_11_), .F3(dummy_abc_12_) );
      defparam ii0885.CONFIG_DATA = 16'hFFFF;
      defparam ii0885.PLACE_LOCATION = "NONE";
      defparam ii0885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0886 ( .DX(nn0886), .F0(xBgn[0]), .F1(xEnd[0]), .F2(dummy_abc_13_), .F3(dummy_abc_14_) );
      defparam ii0886.CONFIG_DATA = 16'h6666;
      defparam ii0886.PLACE_LOCATION = "NONE";
      defparam ii0886.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0887 ( .DX(nn0887), .F0(\cal1_v__reg[11]|Q_net ), .F1(nn0886), .F2(dummy_abc_15_), .F3(dummy_abc_16_) );
      defparam ii0887.CONFIG_DATA = 16'h6666;
      defparam ii0887.PLACE_LOCATION = "NONE";
      defparam ii0887.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0888 ( .DX(nn0888), .F0(nn0886), .F1(dummy_abc_17_), .F2(dummy_abc_18_), .F3(dummy_abc_19_) );
      defparam ii0888.CONFIG_DATA = 16'h5555;
      defparam ii0888.PLACE_LOCATION = "NONE";
      defparam ii0888.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0889 ( .DX(nn0889), .F0(xBgn[1]), .F1(xEnd[1]), .F2(dummy_abc_20_), .F3(dummy_abc_21_) );
      defparam ii0889.CONFIG_DATA = 16'h9999;
      defparam ii0889.PLACE_LOCATION = "NONE";
      defparam ii0889.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0890 ( .DX(nn0890), .F0(xBgn[2]), .F1(xEnd[2]), .F2(dummy_abc_22_), .F3(dummy_abc_23_) );
      defparam ii0890.CONFIG_DATA = 16'h9999;
      defparam ii0890.PLACE_LOCATION = "NONE";
      defparam ii0890.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0891 ( .DX(nn0891), .F0(xBgn[3]), .F1(xEnd[3]), .F2(dummy_abc_24_), .F3(dummy_abc_25_) );
      defparam ii0891.CONFIG_DATA = 16'h9999;
      defparam ii0891.PLACE_LOCATION = "NONE";
      defparam ii0891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0892 ( .DX(nn0892), .F0(xBgn[4]), .F1(xEnd[4]), .F2(dummy_abc_26_), .F3(dummy_abc_27_) );
      defparam ii0892.CONFIG_DATA = 16'h9999;
      defparam ii0892.PLACE_LOCATION = "NONE";
      defparam ii0892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0893 ( .DX(nn0893), .F0(xBgn[5]), .F1(xEnd[5]), .F2(dummy_abc_28_), .F3(dummy_abc_29_) );
      defparam ii0893.CONFIG_DATA = 16'h9999;
      defparam ii0893.PLACE_LOCATION = "NONE";
      defparam ii0893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0894 ( .DX(nn0894), .F0(xBgn[6]), .F1(xEnd[6]), .F2(dummy_abc_30_), .F3(dummy_abc_31_) );
      defparam ii0894.CONFIG_DATA = 16'h9999;
      defparam ii0894.PLACE_LOCATION = "NONE";
      defparam ii0894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0895 ( .DX(nn0895), .F0(xBgn[7]), .F1(xEnd[7]), .F2(dummy_abc_32_), .F3(dummy_abc_33_) );
      defparam ii0895.CONFIG_DATA = 16'h9999;
      defparam ii0895.PLACE_LOCATION = "NONE";
      defparam ii0895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0896 ( .DX(nn0896), .F0(xBgn[8]), .F1(xEnd[8]), .F2(dummy_abc_34_), .F3(dummy_abc_35_) );
      defparam ii0896.CONFIG_DATA = 16'h9999;
      defparam ii0896.PLACE_LOCATION = "NONE";
      defparam ii0896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0897 ( .DX(nn0897), .F0(xBgn[9]), .F1(xEnd[9]), .F2(dummy_abc_36_), .F3(dummy_abc_37_) );
      defparam ii0897.CONFIG_DATA = 16'h9999;
      defparam ii0897.PLACE_LOCATION = "NONE";
      defparam ii0897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0898 ( .DX(nn0898), .F0(xBgn[10]), .F1(xEnd[10]), .F2(dummy_abc_38_), .F3(dummy_abc_39_) );
      defparam ii0898.CONFIG_DATA = 16'h9999;
      defparam ii0898.PLACE_LOCATION = "NONE";
      defparam ii0898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0899 ( .DX(nn0899), .F0(dummy_abc_40_), .F1(dummy_abc_41_), .F2(dummy_abc_42_), .F3(dummy_abc_43_) );
      defparam ii0899.CONFIG_DATA = 16'hFFFF;
      defparam ii0899.PLACE_LOCATION = "NONE";
      defparam ii0899.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_293_ ( 
        .CA( {a_acc_en_cal1_u137_mac, xEnd[10], xEnd[9], xEnd[8], xEnd[7], 
              xEnd[6], xEnd[5], xEnd[4], xEnd[3], xEnd[2], xEnd[1], xEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_133_ ), 
        .DX( {nn0899, nn0898, nn0897, nn0896, nn0895, nn0894, nn0893, nn0892, 
              nn0891, nn0890, nn0889, nn0888} ), 
        .SUM( {\u2_XORCI_11|SUM_net , \u2_XORCI_10|SUM_net , \u2_XORCI_9|SUM_net , 
              \u2_XORCI_8|SUM_net , \u2_XORCI_7|SUM_net , \u2_XORCI_6|SUM_net , 
              \u2_XORCI_5|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_3|SUM_net , 
              \u2_XORCI_2|SUM_net , \u2_XORCI_1|SUM_net , \u2_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0914 ( .DX(nn0914), .F0(xBgn[0]), .F1(xEnd[0]), .F2(dummy_abc_44_), .F3(dummy_abc_45_) );
      defparam ii0914.CONFIG_DATA = 16'h6666;
      defparam ii0914.PLACE_LOCATION = "NONE";
      defparam ii0914.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0915 ( .DX(nn0915), .F0(\u2_XORCI_1|SUM_net ), .F1(dummy_abc_46_), .F2(dummy_abc_47_), .F3(dummy_abc_48_) );
      defparam ii0915.CONFIG_DATA = 16'h5555;
      defparam ii0915.PLACE_LOCATION = "NONE";
      defparam ii0915.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0916 ( .DX(nn0916), .F0(\u2_XORCI_2|SUM_net ), .F1(dummy_abc_49_), .F2(dummy_abc_50_), .F3(dummy_abc_51_) );
      defparam ii0916.CONFIG_DATA = 16'h5555;
      defparam ii0916.PLACE_LOCATION = "NONE";
      defparam ii0916.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0917 ( .DX(nn0917), .F0(\u2_XORCI_3|SUM_net ), .F1(dummy_abc_52_), .F2(dummy_abc_53_), .F3(dummy_abc_54_) );
      defparam ii0917.CONFIG_DATA = 16'h5555;
      defparam ii0917.PLACE_LOCATION = "NONE";
      defparam ii0917.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0918 ( .DX(nn0918), .F0(\u2_XORCI_4|SUM_net ), .F1(dummy_abc_55_), .F2(dummy_abc_56_), .F3(dummy_abc_57_) );
      defparam ii0918.CONFIG_DATA = 16'h5555;
      defparam ii0918.PLACE_LOCATION = "NONE";
      defparam ii0918.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0919 ( .DX(nn0919), .F0(\u2_XORCI_5|SUM_net ), .F1(dummy_abc_58_), .F2(dummy_abc_59_), .F3(dummy_abc_60_) );
      defparam ii0919.CONFIG_DATA = 16'h5555;
      defparam ii0919.PLACE_LOCATION = "NONE";
      defparam ii0919.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0920 ( .DX(nn0920), .F0(\u2_XORCI_6|SUM_net ), .F1(dummy_abc_61_), .F2(dummy_abc_62_), .F3(dummy_abc_63_) );
      defparam ii0920.CONFIG_DATA = 16'h5555;
      defparam ii0920.PLACE_LOCATION = "NONE";
      defparam ii0920.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0921 ( .DX(nn0921), .F0(\u2_XORCI_7|SUM_net ), .F1(dummy_abc_64_), .F2(dummy_abc_65_), .F3(dummy_abc_66_) );
      defparam ii0921.CONFIG_DATA = 16'h5555;
      defparam ii0921.PLACE_LOCATION = "NONE";
      defparam ii0921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0922 ( .DX(nn0922), .F0(\u2_XORCI_8|SUM_net ), .F1(dummy_abc_67_), .F2(dummy_abc_68_), .F3(dummy_abc_69_) );
      defparam ii0922.CONFIG_DATA = 16'h5555;
      defparam ii0922.PLACE_LOCATION = "NONE";
      defparam ii0922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0923 ( .DX(nn0923), .F0(\u2_XORCI_9|SUM_net ), .F1(dummy_abc_70_), .F2(dummy_abc_71_), .F3(dummy_abc_72_) );
      defparam ii0923.CONFIG_DATA = 16'h5555;
      defparam ii0923.PLACE_LOCATION = "NONE";
      defparam ii0923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0924 ( .DX(nn0924), .F0(\u2_XORCI_10|SUM_net ), .F1(dummy_abc_73_), .F2(dummy_abc_74_), .F3(dummy_abc_75_) );
      defparam ii0924.CONFIG_DATA = 16'h5555;
      defparam ii0924.PLACE_LOCATION = "NONE";
      defparam ii0924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0925 ( .DX(nn0925), .F0(dummy_abc_76_), .F1(dummy_abc_77_), .F2(dummy_abc_78_), .F3(dummy_abc_79_) );
      defparam ii0925.CONFIG_DATA = 16'h0000;
      defparam ii0925.PLACE_LOCATION = "NONE";
      defparam ii0925.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_294_ ( 
        .CA( {\u2_XORCI_11|SUM_net , \u2_XORCI_10|SUM_net , \u2_XORCI_9|SUM_net , 
              \u2_XORCI_8|SUM_net , \u2_XORCI_7|SUM_net , \u2_XORCI_6|SUM_net , 
              \u2_XORCI_5|SUM_net , \u2_XORCI_4|SUM_net , \u2_XORCI_3|SUM_net , 
              \u2_XORCI_2|SUM_net , \u2_XORCI_1|SUM_net , nn0886} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_134_ ), 
        .DX( {nn0925, nn0924, nn0923, nn0922, nn0921, nn0920, nn0919, nn0918, 
              nn0917, nn0916, nn0915, nn0914} ), 
        .SUM( {dummy_135_, \u3_XORCI_10|SUM_net , \u3_XORCI_9|SUM_net , 
              \u3_XORCI_8|SUM_net , \u3_XORCI_7|SUM_net , \u3_XORCI_6|SUM_net , 
              \u3_XORCI_5|SUM_net , \u3_XORCI_4|SUM_net , \u3_XORCI_3|SUM_net , 
              \u3_XORCI_2|SUM_net , \u3_XORCI_1|SUM_net , \u3_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii0940 ( .DX(nn0940), .F0(\cal1_v__reg[12]|Q_net ), .F1(\u3_XORCI_1|SUM_net ), .F2(dummy_abc_80_), .F3(dummy_abc_81_) );
      defparam ii0940.CONFIG_DATA = 16'h9999;
      defparam ii0940.PLACE_LOCATION = "NONE";
      defparam ii0940.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0941 ( .DX(nn0941), .F0(\cal1_v__reg[13]|Q_net ), .F1(\u3_XORCI_2|SUM_net ), .F2(dummy_abc_82_), .F3(dummy_abc_83_) );
      defparam ii0941.CONFIG_DATA = 16'h9999;
      defparam ii0941.PLACE_LOCATION = "NONE";
      defparam ii0941.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0942 ( .DX(nn0942), .F0(\cal1_v__reg[14]|Q_net ), .F1(\u3_XORCI_3|SUM_net ), .F2(dummy_abc_84_), .F3(dummy_abc_85_) );
      defparam ii0942.CONFIG_DATA = 16'h9999;
      defparam ii0942.PLACE_LOCATION = "NONE";
      defparam ii0942.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0943 ( .DX(nn0943), .F0(\cal1_v__reg[15]|Q_net ), .F1(\u3_XORCI_4|SUM_net ), .F2(dummy_abc_86_), .F3(dummy_abc_87_) );
      defparam ii0943.CONFIG_DATA = 16'h9999;
      defparam ii0943.PLACE_LOCATION = "NONE";
      defparam ii0943.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0944 ( .DX(nn0944), .F0(\cal1_v__reg[16]|Q_net ), .F1(\u3_XORCI_5|SUM_net ), .F2(dummy_abc_88_), .F3(dummy_abc_89_) );
      defparam ii0944.CONFIG_DATA = 16'h9999;
      defparam ii0944.PLACE_LOCATION = "NONE";
      defparam ii0944.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0945 ( .DX(nn0945), .F0(\u3_XORCI_6|SUM_net ), .F1(dummy_abc_90_), .F2(dummy_abc_91_), .F3(dummy_abc_92_) );
      defparam ii0945.CONFIG_DATA = 16'h5555;
      defparam ii0945.PLACE_LOCATION = "NONE";
      defparam ii0945.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0946 ( .DX(nn0946), .F0(\u3_XORCI_7|SUM_net ), .F1(dummy_abc_93_), .F2(dummy_abc_94_), .F3(dummy_abc_95_) );
      defparam ii0946.CONFIG_DATA = 16'h5555;
      defparam ii0946.PLACE_LOCATION = "NONE";
      defparam ii0946.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0947 ( .DX(nn0947), .F0(\u3_XORCI_8|SUM_net ), .F1(dummy_abc_96_), .F2(dummy_abc_97_), .F3(dummy_abc_98_) );
      defparam ii0947.CONFIG_DATA = 16'h5555;
      defparam ii0947.PLACE_LOCATION = "NONE";
      defparam ii0947.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0948 ( .DX(nn0948), .F0(\u3_XORCI_9|SUM_net ), .F1(dummy_abc_99_), .F2(dummy_abc_100_), .F3(dummy_abc_101_) );
      defparam ii0948.CONFIG_DATA = 16'h5555;
      defparam ii0948.PLACE_LOCATION = "NONE";
      defparam ii0948.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0949 ( .DX(nn0949), .F0(\u3_XORCI_10|SUM_net ), .F1(dummy_abc_102_), .F2(dummy_abc_103_), .F3(dummy_abc_104_) );
      defparam ii0949.CONFIG_DATA = 16'h5555;
      defparam ii0949.PLACE_LOCATION = "NONE";
      defparam ii0949.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0950 ( .DX(nn0950), .F0(dummy_abc_105_), .F1(dummy_abc_106_), .F2(dummy_abc_107_), .F3(dummy_abc_108_) );
      defparam ii0950.CONFIG_DATA = 16'hFFFF;
      defparam ii0950.PLACE_LOCATION = "NONE";
      defparam ii0950.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_213_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, \cal1_v__reg[16]|Q_net , \cal1_v__reg[15]|Q_net , 
              \cal1_v__reg[14]|Q_net , \cal1_v__reg[13]|Q_net , \cal1_v__reg[12]|Q_net , 
              \cal1_v__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_62_ ), 
        .DX( {nn0950, nn0949, nn0948, nn0947, nn0946, nn0945, nn0944, nn0943, 
              nn0942, nn0941, nn0940, nn0887} ), 
        .SUM( {\cal1_u63_XORCI_11|SUM_net , dummy_63_, dummy_64_, dummy_65_, 
              dummy_66_, dummy_67_, dummy_68_, dummy_69_, dummy_70_, dummy_71_, 
              dummy_72_, dummy_73_} )
      );
    CS_LUT4_PRIM ii0965 ( .DX(nn0965), .F0(\c1r2_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_109_) );
      defparam ii0965.CONFIG_DATA = 16'hCACA;
      defparam ii0965.PLACE_LOCATION = "NONE";
      defparam ii0965.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0966 ( .DX(\a_dinx[0]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u138_mac ), .F3(nn0965) );
      defparam ii0966.CONFIG_DATA = 16'hE4A0;
      defparam ii0966.PLACE_LOCATION = "NONE";
      defparam ii0966.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0967 ( .DX(nn0967), .F0(\c1r2_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_110_) );
      defparam ii0967.CONFIG_DATA = 16'hCACA;
      defparam ii0967.PLACE_LOCATION = "NONE";
      defparam ii0967.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0968 ( .DX(\a_dinx[0]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u139_mac ), .F3(nn0967) );
      defparam ii0968.CONFIG_DATA = 16'hE4A0;
      defparam ii0968.PLACE_LOCATION = "NONE";
      defparam ii0968.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0969 ( .DX(\a_dinx[0]_cal1_u142_mac ), .F0(\c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0969.CONFIG_DATA = 16'hCA00;
      defparam ii0969.PLACE_LOCATION = "NONE";
      defparam ii0969.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0970 ( .DX(\a_dinx[0]_cal1_u143_mac ), .F0(\c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0970.CONFIG_DATA = 16'hCA00;
      defparam ii0970.PLACE_LOCATION = "NONE";
      defparam ii0970.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0971 ( .DX(nn0971), .F0(\c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_111_) );
      defparam ii0971.CONFIG_DATA = 16'hCACA;
      defparam ii0971.PLACE_LOCATION = "NONE";
      defparam ii0971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0972 ( .DX(\a_dinx[0]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u142_mac ), .F3(nn0971) );
      defparam ii0972.CONFIG_DATA = 16'hE4A0;
      defparam ii0972.PLACE_LOCATION = "NONE";
      defparam ii0972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0973 ( .DX(nn0973), .F0(\c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_112_) );
      defparam ii0973.CONFIG_DATA = 16'hCACA;
      defparam ii0973.PLACE_LOCATION = "NONE";
      defparam ii0973.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0974 ( .DX(\a_dinx[0]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u143_mac ), .F3(nn0973) );
      defparam ii0974.CONFIG_DATA = 16'hE4A0;
      defparam ii0974.PLACE_LOCATION = "NONE";
      defparam ii0974.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0975 ( .DX(\a_dinx[0]_cal1_u146_mac ), .F0(\c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0975.CONFIG_DATA = 16'hCA00;
      defparam ii0975.PLACE_LOCATION = "NONE";
      defparam ii0975.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0976 ( .DX(\a_dinx[0]_cal1_u147_mac ), .F0(\c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0976.CONFIG_DATA = 16'hCA00;
      defparam ii0976.PLACE_LOCATION = "NONE";
      defparam ii0976.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0977 ( .DX(nn0977), .F0(\c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_113_) );
      defparam ii0977.CONFIG_DATA = 16'hCACA;
      defparam ii0977.PLACE_LOCATION = "NONE";
      defparam ii0977.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0978 ( .DX(\a_dinx[0]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u146_mac ), .F3(nn0977) );
      defparam ii0978.CONFIG_DATA = 16'hE4A0;
      defparam ii0978.PLACE_LOCATION = "NONE";
      defparam ii0978.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0979 ( .DX(nn0979), .F0(\c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_114_) );
      defparam ii0979.CONFIG_DATA = 16'hCACA;
      defparam ii0979.PLACE_LOCATION = "NONE";
      defparam ii0979.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0980 ( .DX(\a_dinx[0]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[0]_cal1_u147_mac ), .F3(nn0979) );
      defparam ii0980.CONFIG_DATA = 16'hE4A0;
      defparam ii0980.PLACE_LOCATION = "NONE";
      defparam ii0980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0981 ( .DX(\a_dinx[1]_cal1_u138_mac ), .F0(\c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0981.CONFIG_DATA = 16'hCA00;
      defparam ii0981.PLACE_LOCATION = "NONE";
      defparam ii0981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0982 ( .DX(\a_dinx[1]_cal1_u139_mac ), .F0(\c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0982.CONFIG_DATA = 16'hCA00;
      defparam ii0982.PLACE_LOCATION = "NONE";
      defparam ii0982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0983 ( .DX(nn0983), .F0(\c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_115_) );
      defparam ii0983.CONFIG_DATA = 16'hCACA;
      defparam ii0983.PLACE_LOCATION = "NONE";
      defparam ii0983.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0984 ( .DX(\a_dinx[1]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u138_mac ), .F3(nn0983) );
      defparam ii0984.CONFIG_DATA = 16'hE4A0;
      defparam ii0984.PLACE_LOCATION = "NONE";
      defparam ii0984.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0985 ( .DX(nn0985), .F0(\c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_116_) );
      defparam ii0985.CONFIG_DATA = 16'hCACA;
      defparam ii0985.PLACE_LOCATION = "NONE";
      defparam ii0985.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0986 ( .DX(\a_dinx[1]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u139_mac ), .F3(nn0985) );
      defparam ii0986.CONFIG_DATA = 16'hE4A0;
      defparam ii0986.PLACE_LOCATION = "NONE";
      defparam ii0986.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0987 ( .DX(\a_dinx[1]_cal1_u142_mac ), .F0(\c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0987.CONFIG_DATA = 16'hCA00;
      defparam ii0987.PLACE_LOCATION = "NONE";
      defparam ii0987.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0988 ( .DX(\a_dinx[1]_cal1_u143_mac ), .F0(\c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0988.CONFIG_DATA = 16'hCA00;
      defparam ii0988.PLACE_LOCATION = "NONE";
      defparam ii0988.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0989 ( .DX(nn0989), .F0(\c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_117_) );
      defparam ii0989.CONFIG_DATA = 16'hCACA;
      defparam ii0989.PLACE_LOCATION = "NONE";
      defparam ii0989.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0990 ( .DX(\a_dinx[1]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u142_mac ), .F3(nn0989) );
      defparam ii0990.CONFIG_DATA = 16'hE4A0;
      defparam ii0990.PLACE_LOCATION = "NONE";
      defparam ii0990.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0991 ( .DX(nn0991), .F0(\c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_118_) );
      defparam ii0991.CONFIG_DATA = 16'hCACA;
      defparam ii0991.PLACE_LOCATION = "NONE";
      defparam ii0991.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0992 ( .DX(\a_dinx[1]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u143_mac ), .F3(nn0991) );
      defparam ii0992.CONFIG_DATA = 16'hE4A0;
      defparam ii0992.PLACE_LOCATION = "NONE";
      defparam ii0992.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0993 ( .DX(\a_dinx[1]_cal1_u146_mac ), .F0(\c1r2_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0993.CONFIG_DATA = 16'hCA00;
      defparam ii0993.PLACE_LOCATION = "NONE";
      defparam ii0993.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0994 ( .DX(\a_dinx[1]_cal1_u147_mac ), .F0(\c1r2_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0994.CONFIG_DATA = 16'hCA00;
      defparam ii0994.PLACE_LOCATION = "NONE";
      defparam ii0994.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0995 ( .DX(nn0995), .F0(\c1r2_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_119_) );
      defparam ii0995.CONFIG_DATA = 16'hCACA;
      defparam ii0995.PLACE_LOCATION = "NONE";
      defparam ii0995.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0996 ( .DX(\a_dinx[1]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u146_mac ), .F3(nn0995) );
      defparam ii0996.CONFIG_DATA = 16'hE4A0;
      defparam ii0996.PLACE_LOCATION = "NONE";
      defparam ii0996.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0997 ( .DX(nn0997), .F0(\c1r2_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_120_) );
      defparam ii0997.CONFIG_DATA = 16'hCACA;
      defparam ii0997.PLACE_LOCATION = "NONE";
      defparam ii0997.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0998 ( .DX(\a_dinx[1]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[1]_cal1_u147_mac ), .F3(nn0997) );
      defparam ii0998.CONFIG_DATA = 16'hE4A0;
      defparam ii0998.PLACE_LOCATION = "NONE";
      defparam ii0998.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii0999 ( .DX(\a_dinx[2]_cal1_u138_mac ), .F0(\c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii0999.CONFIG_DATA = 16'hCA00;
      defparam ii0999.PLACE_LOCATION = "NONE";
      defparam ii0999.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1000 ( .DX(\a_dinx[2]_cal1_u139_mac ), .F0(\c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1000.CONFIG_DATA = 16'hCA00;
      defparam ii1000.PLACE_LOCATION = "NONE";
      defparam ii1000.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1001 ( .DX(nn1001), .F0(\c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_121_) );
      defparam ii1001.CONFIG_DATA = 16'hCACA;
      defparam ii1001.PLACE_LOCATION = "NONE";
      defparam ii1001.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1002 ( .DX(\a_dinx[2]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u138_mac ), .F3(nn1001) );
      defparam ii1002.CONFIG_DATA = 16'hE4A0;
      defparam ii1002.PLACE_LOCATION = "NONE";
      defparam ii1002.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1003 ( .DX(nn1003), .F0(\c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_122_) );
      defparam ii1003.CONFIG_DATA = 16'hCACA;
      defparam ii1003.PLACE_LOCATION = "NONE";
      defparam ii1003.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1004 ( .DX(\a_dinx[2]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u139_mac ), .F3(nn1003) );
      defparam ii1004.CONFIG_DATA = 16'hE4A0;
      defparam ii1004.PLACE_LOCATION = "NONE";
      defparam ii1004.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1005 ( .DX(\a_dinx[2]_cal1_u142_mac ), .F0(\c1r2_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1005.CONFIG_DATA = 16'hCA00;
      defparam ii1005.PLACE_LOCATION = "NONE";
      defparam ii1005.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1006 ( .DX(\a_dinx[2]_cal1_u143_mac ), .F0(\c1r2_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1006.CONFIG_DATA = 16'hCA00;
      defparam ii1006.PLACE_LOCATION = "NONE";
      defparam ii1006.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1007 ( .DX(nn1007), .F0(\c1r2_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_123_) );
      defparam ii1007.CONFIG_DATA = 16'hCACA;
      defparam ii1007.PLACE_LOCATION = "NONE";
      defparam ii1007.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1008 ( .DX(\a_dinx[2]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u142_mac ), .F3(nn1007) );
      defparam ii1008.CONFIG_DATA = 16'hE4A0;
      defparam ii1008.PLACE_LOCATION = "NONE";
      defparam ii1008.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1009 ( .DX(nn1009), .F0(\c1r2_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_124_) );
      defparam ii1009.CONFIG_DATA = 16'hCACA;
      defparam ii1009.PLACE_LOCATION = "NONE";
      defparam ii1009.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1010 ( .DX(\a_dinx[2]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u143_mac ), .F3(nn1009) );
      defparam ii1010.CONFIG_DATA = 16'hE4A0;
      defparam ii1010.PLACE_LOCATION = "NONE";
      defparam ii1010.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1011 ( .DX(\a_dinx[2]_cal1_u146_mac ), .F0(\c1r1_q[0]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1011.CONFIG_DATA = 16'hCA00;
      defparam ii1011.PLACE_LOCATION = "NONE";
      defparam ii1011.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1012 ( .DX(\a_dinx[2]_cal1_u147_mac ), .F0(\c1r1_q[9]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1012.CONFIG_DATA = 16'hCA00;
      defparam ii1012.PLACE_LOCATION = "NONE";
      defparam ii1012.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1013 ( .DX(nn1013), .F0(\c1r1_q[0]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_125_) );
      defparam ii1013.CONFIG_DATA = 16'hCACA;
      defparam ii1013.PLACE_LOCATION = "NONE";
      defparam ii1013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1014 ( .DX(\a_dinx[2]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u146_mac ), .F3(nn1013) );
      defparam ii1014.CONFIG_DATA = 16'hE4A0;
      defparam ii1014.PLACE_LOCATION = "NONE";
      defparam ii1014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1015 ( .DX(nn1015), .F0(\c1r1_q[9]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_126_) );
      defparam ii1015.CONFIG_DATA = 16'hCACA;
      defparam ii1015.PLACE_LOCATION = "NONE";
      defparam ii1015.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1016 ( .DX(\a_dinx[2]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[2]_cal1_u147_mac ), .F3(nn1015) );
      defparam ii1016.CONFIG_DATA = 16'hE4A0;
      defparam ii1016.PLACE_LOCATION = "NONE";
      defparam ii1016.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1017 ( .DX(\a_dinx[3]_cal1_u138_mac ), .F0(\c1r2_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1017.CONFIG_DATA = 16'hCA00;
      defparam ii1017.PLACE_LOCATION = "NONE";
      defparam ii1017.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1018 ( .DX(\a_dinx[3]_cal1_u139_mac ), .F0(\c1r2_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1018.CONFIG_DATA = 16'hCA00;
      defparam ii1018.PLACE_LOCATION = "NONE";
      defparam ii1018.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1019 ( .DX(nn1019), .F0(\c1r2_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_127_) );
      defparam ii1019.CONFIG_DATA = 16'hCACA;
      defparam ii1019.PLACE_LOCATION = "NONE";
      defparam ii1019.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1020 ( .DX(\a_dinx[3]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u138_mac ), .F3(nn1019) );
      defparam ii1020.CONFIG_DATA = 16'hE4A0;
      defparam ii1020.PLACE_LOCATION = "NONE";
      defparam ii1020.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1021 ( .DX(nn1021), .F0(\c1r2_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_128_) );
      defparam ii1021.CONFIG_DATA = 16'hCACA;
      defparam ii1021.PLACE_LOCATION = "NONE";
      defparam ii1021.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1022 ( .DX(\a_dinx[3]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u139_mac ), .F3(nn1021) );
      defparam ii1022.CONFIG_DATA = 16'hE4A0;
      defparam ii1022.PLACE_LOCATION = "NONE";
      defparam ii1022.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1023 ( .DX(\a_dinx[3]_cal1_u142_mac ), .F0(\c1r1_q[3]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1023.CONFIG_DATA = 16'hCA00;
      defparam ii1023.PLACE_LOCATION = "NONE";
      defparam ii1023.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1024 ( .DX(\a_dinx[3]_cal1_u143_mac ), .F0(\c1r1_q[12]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1024.CONFIG_DATA = 16'hCA00;
      defparam ii1024.PLACE_LOCATION = "NONE";
      defparam ii1024.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1025 ( .DX(nn1025), .F0(\c1r1_q[3]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_129_) );
      defparam ii1025.CONFIG_DATA = 16'hCACA;
      defparam ii1025.PLACE_LOCATION = "NONE";
      defparam ii1025.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1026 ( .DX(\a_dinx[3]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u142_mac ), .F3(nn1025) );
      defparam ii1026.CONFIG_DATA = 16'hE4A0;
      defparam ii1026.PLACE_LOCATION = "NONE";
      defparam ii1026.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1027 ( .DX(nn1027), .F0(\c1r1_q[12]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_130_) );
      defparam ii1027.CONFIG_DATA = 16'hCACA;
      defparam ii1027.PLACE_LOCATION = "NONE";
      defparam ii1027.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1028 ( .DX(\a_dinx[3]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u143_mac ), .F3(nn1027) );
      defparam ii1028.CONFIG_DATA = 16'hE4A0;
      defparam ii1028.PLACE_LOCATION = "NONE";
      defparam ii1028.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1029 ( .DX(\a_dinx[3]_cal1_u146_mac ), .F0(\c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1029.CONFIG_DATA = 16'hCA00;
      defparam ii1029.PLACE_LOCATION = "NONE";
      defparam ii1029.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1030 ( .DX(\a_dinx[3]_cal1_u147_mac ), .F0(\c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1030.CONFIG_DATA = 16'hCA00;
      defparam ii1030.PLACE_LOCATION = "NONE";
      defparam ii1030.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1031 ( .DX(nn1031), .F0(\c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_131_) );
      defparam ii1031.CONFIG_DATA = 16'hCACA;
      defparam ii1031.PLACE_LOCATION = "NONE";
      defparam ii1031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1032 ( .DX(\a_dinx[3]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u146_mac ), .F3(nn1031) );
      defparam ii1032.CONFIG_DATA = 16'hE4A0;
      defparam ii1032.PLACE_LOCATION = "NONE";
      defparam ii1032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1033 ( .DX(nn1033), .F0(\c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_132_) );
      defparam ii1033.CONFIG_DATA = 16'hCACA;
      defparam ii1033.PLACE_LOCATION = "NONE";
      defparam ii1033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1034 ( .DX(\a_dinx[3]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[3]_cal1_u147_mac ), .F3(nn1033) );
      defparam ii1034.CONFIG_DATA = 16'hE4A0;
      defparam ii1034.PLACE_LOCATION = "NONE";
      defparam ii1034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1035 ( .DX(\a_dinx[4]_cal1_u138_mac ), .F0(\c1r1_q[2]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1035.CONFIG_DATA = 16'hCA00;
      defparam ii1035.PLACE_LOCATION = "NONE";
      defparam ii1035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1036 ( .DX(\a_dinx[4]_cal1_u139_mac ), .F0(\c1r1_q[11]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1036.CONFIG_DATA = 16'hCA00;
      defparam ii1036.PLACE_LOCATION = "NONE";
      defparam ii1036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1037 ( .DX(nn1037), .F0(\c1r1_q[2]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_133_) );
      defparam ii1037.CONFIG_DATA = 16'hCACA;
      defparam ii1037.PLACE_LOCATION = "NONE";
      defparam ii1037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1038 ( .DX(\a_dinx[4]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u138_mac ), .F3(nn1037) );
      defparam ii1038.CONFIG_DATA = 16'hE4A0;
      defparam ii1038.PLACE_LOCATION = "NONE";
      defparam ii1038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1039 ( .DX(nn1039), .F0(\c1r1_q[11]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_134_) );
      defparam ii1039.CONFIG_DATA = 16'hCACA;
      defparam ii1039.PLACE_LOCATION = "NONE";
      defparam ii1039.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1040 ( .DX(\a_dinx[4]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u139_mac ), .F3(nn1039) );
      defparam ii1040.CONFIG_DATA = 16'hE4A0;
      defparam ii1040.PLACE_LOCATION = "NONE";
      defparam ii1040.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1041 ( .DX(\a_dinx[4]_cal1_u142_mac ), .F0(\c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1041.CONFIG_DATA = 16'hCA00;
      defparam ii1041.PLACE_LOCATION = "NONE";
      defparam ii1041.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1042 ( .DX(\a_dinx[4]_cal1_u143_mac ), .F0(\c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1042.CONFIG_DATA = 16'hCA00;
      defparam ii1042.PLACE_LOCATION = "NONE";
      defparam ii1042.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1043 ( .DX(nn1043), .F0(\c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_135_) );
      defparam ii1043.CONFIG_DATA = 16'hCACA;
      defparam ii1043.PLACE_LOCATION = "NONE";
      defparam ii1043.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1044 ( .DX(\a_dinx[4]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u142_mac ), .F3(nn1043) );
      defparam ii1044.CONFIG_DATA = 16'hE4A0;
      defparam ii1044.PLACE_LOCATION = "NONE";
      defparam ii1044.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1045 ( .DX(nn1045), .F0(\c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_136_) );
      defparam ii1045.CONFIG_DATA = 16'hCACA;
      defparam ii1045.PLACE_LOCATION = "NONE";
      defparam ii1045.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1046 ( .DX(\a_dinx[4]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u143_mac ), .F3(nn1045) );
      defparam ii1046.CONFIG_DATA = 16'hE4A0;
      defparam ii1046.PLACE_LOCATION = "NONE";
      defparam ii1046.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1047 ( .DX(\a_dinx[4]_cal1_u146_mac ), .F0(\c1r2_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1047.CONFIG_DATA = 16'hCA00;
      defparam ii1047.PLACE_LOCATION = "NONE";
      defparam ii1047.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1048 ( .DX(\a_dinx[4]_cal1_u147_mac ), .F0(\c1r2_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1048.CONFIG_DATA = 16'hCA00;
      defparam ii1048.PLACE_LOCATION = "NONE";
      defparam ii1048.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1049 ( .DX(nn1049), .F0(\c1r2_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[1]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_137_) );
      defparam ii1049.CONFIG_DATA = 16'hCACA;
      defparam ii1049.PLACE_LOCATION = "NONE";
      defparam ii1049.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1050 ( .DX(\a_dinx[4]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u146_mac ), .F3(nn1049) );
      defparam ii1050.CONFIG_DATA = 16'hE4A0;
      defparam ii1050.PLACE_LOCATION = "NONE";
      defparam ii1050.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1051 ( .DX(nn1051), .F0(\c1r2_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[10]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_138_) );
      defparam ii1051.CONFIG_DATA = 16'hCACA;
      defparam ii1051.PLACE_LOCATION = "NONE";
      defparam ii1051.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1052 ( .DX(\a_dinx[4]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[4]_cal1_u147_mac ), .F3(nn1051) );
      defparam ii1052.CONFIG_DATA = 16'hE4A0;
      defparam ii1052.PLACE_LOCATION = "NONE";
      defparam ii1052.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1053 ( .DX(\a_dinx[5]_cal1_u138_mac ), .F0(\c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1053.CONFIG_DATA = 16'hCA00;
      defparam ii1053.PLACE_LOCATION = "NONE";
      defparam ii1053.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1054 ( .DX(\a_dinx[5]_cal1_u139_mac ), .F0(\c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1054.CONFIG_DATA = 16'hCA00;
      defparam ii1054.PLACE_LOCATION = "NONE";
      defparam ii1054.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1055 ( .DX(nn1055), .F0(\c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_139_) );
      defparam ii1055.CONFIG_DATA = 16'hCACA;
      defparam ii1055.PLACE_LOCATION = "NONE";
      defparam ii1055.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1056 ( .DX(\a_dinx[5]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u138_mac ), .F3(nn1055) );
      defparam ii1056.CONFIG_DATA = 16'hE4A0;
      defparam ii1056.PLACE_LOCATION = "NONE";
      defparam ii1056.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1057 ( .DX(nn1057), .F0(\c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_140_) );
      defparam ii1057.CONFIG_DATA = 16'hCACA;
      defparam ii1057.PLACE_LOCATION = "NONE";
      defparam ii1057.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1058 ( .DX(\a_dinx[5]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u139_mac ), .F3(nn1057) );
      defparam ii1058.CONFIG_DATA = 16'hE4A0;
      defparam ii1058.PLACE_LOCATION = "NONE";
      defparam ii1058.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1059 ( .DX(\a_dinx[5]_cal1_u142_mac ), .F0(\c1r2_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1059.CONFIG_DATA = 16'hCA00;
      defparam ii1059.PLACE_LOCATION = "NONE";
      defparam ii1059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1060 ( .DX(\a_dinx[5]_cal1_u143_mac ), .F0(\c1r2_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1060.CONFIG_DATA = 16'hCA00;
      defparam ii1060.PLACE_LOCATION = "NONE";
      defparam ii1060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1061 ( .DX(nn1061), .F0(\c1r2_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[0]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_141_) );
      defparam ii1061.CONFIG_DATA = 16'hCACA;
      defparam ii1061.PLACE_LOCATION = "NONE";
      defparam ii1061.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1062 ( .DX(\a_dinx[5]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u142_mac ), .F3(nn1061) );
      defparam ii1062.CONFIG_DATA = 16'hE4A0;
      defparam ii1062.PLACE_LOCATION = "NONE";
      defparam ii1062.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1063 ( .DX(nn1063), .F0(\c1r2_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[9]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_142_) );
      defparam ii1063.CONFIG_DATA = 16'hCACA;
      defparam ii1063.PLACE_LOCATION = "NONE";
      defparam ii1063.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1064 ( .DX(\a_dinx[5]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u143_mac ), .F3(nn1063) );
      defparam ii1064.CONFIG_DATA = 16'hE4A0;
      defparam ii1064.PLACE_LOCATION = "NONE";
      defparam ii1064.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1065 ( .DX(\a_dinx[5]_cal1_u146_mac ), .F0(\c1r1_q[1]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1065.CONFIG_DATA = 16'hCA00;
      defparam ii1065.PLACE_LOCATION = "NONE";
      defparam ii1065.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1066 ( .DX(\a_dinx[5]_cal1_u147_mac ), .F0(\c1r1_q[10]_fifo1_ram_inst_0B_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0B_u_emb18k_1 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1066.CONFIG_DATA = 16'hCA00;
      defparam ii1066.PLACE_LOCATION = "NONE";
      defparam ii1066.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1067 ( .DX(nn1067), .F0(\c1r1_q[1]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[1]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_143_) );
      defparam ii1067.CONFIG_DATA = 16'hCACA;
      defparam ii1067.PLACE_LOCATION = "NONE";
      defparam ii1067.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1068 ( .DX(\a_dinx[5]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u146_mac ), .F3(nn1067) );
      defparam ii1068.CONFIG_DATA = 16'hE4A0;
      defparam ii1068.PLACE_LOCATION = "NONE";
      defparam ii1068.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1069 ( .DX(nn1069), .F0(\c1r1_q[10]_fifo1_ram_inst_1B_u_emb18k_1 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1B_u_emb18k_1 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_144_) );
      defparam ii1069.CONFIG_DATA = 16'hCACA;
      defparam ii1069.PLACE_LOCATION = "NONE";
      defparam ii1069.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1070 ( .DX(\a_dinx[5]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[5]_cal1_u147_mac ), .F3(nn1069) );
      defparam ii1070.CONFIG_DATA = 16'hE4A0;
      defparam ii1070.PLACE_LOCATION = "NONE";
      defparam ii1070.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1071 ( .DX(\a_dinx[6]_cal1_u138_mac ), .F0(\c1r2_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1071.CONFIG_DATA = 16'hCA00;
      defparam ii1071.PLACE_LOCATION = "NONE";
      defparam ii1071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1072 ( .DX(\a_dinx[6]_cal1_u139_mac ), .F0(\c1r2_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1072.CONFIG_DATA = 16'hCA00;
      defparam ii1072.PLACE_LOCATION = "NONE";
      defparam ii1072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1073 ( .DX(nn1073), .F0(\c1r2_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[3]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_145_) );
      defparam ii1073.CONFIG_DATA = 16'hCACA;
      defparam ii1073.PLACE_LOCATION = "NONE";
      defparam ii1073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1074 ( .DX(\a_dinx[6]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u138_mac ), .F3(nn1073) );
      defparam ii1074.CONFIG_DATA = 16'hE4A0;
      defparam ii1074.PLACE_LOCATION = "NONE";
      defparam ii1074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1075 ( .DX(nn1075), .F0(\c1r2_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r4_q[12]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_146_) );
      defparam ii1075.CONFIG_DATA = 16'hCACA;
      defparam ii1075.PLACE_LOCATION = "NONE";
      defparam ii1075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1076 ( .DX(\a_dinx[6]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u139_mac ), .F3(nn1075) );
      defparam ii1076.CONFIG_DATA = 16'hE4A0;
      defparam ii1076.PLACE_LOCATION = "NONE";
      defparam ii1076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1077 ( .DX(\a_dinx[6]_cal1_u142_mac ), .F0(\c1r1_q[0]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1077.CONFIG_DATA = 16'hCA00;
      defparam ii1077.PLACE_LOCATION = "NONE";
      defparam ii1077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1078 ( .DX(\a_dinx[6]_cal1_u143_mac ), .F0(\c1r1_q[9]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1078.CONFIG_DATA = 16'hCA00;
      defparam ii1078.PLACE_LOCATION = "NONE";
      defparam ii1078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1079 ( .DX(nn1079), .F0(\c1r1_q[0]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[0]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_147_) );
      defparam ii1079.CONFIG_DATA = 16'hCACA;
      defparam ii1079.PLACE_LOCATION = "NONE";
      defparam ii1079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1080 ( .DX(\a_dinx[6]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u142_mac ), .F3(nn1079) );
      defparam ii1080.CONFIG_DATA = 16'hE4A0;
      defparam ii1080.PLACE_LOCATION = "NONE";
      defparam ii1080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1081 ( .DX(nn1081), .F0(\c1r1_q[9]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[9]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_148_) );
      defparam ii1081.CONFIG_DATA = 16'hCACA;
      defparam ii1081.PLACE_LOCATION = "NONE";
      defparam ii1081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1082 ( .DX(\a_dinx[6]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u143_mac ), .F3(nn1081) );
      defparam ii1082.CONFIG_DATA = 16'hE4A0;
      defparam ii1082.PLACE_LOCATION = "NONE";
      defparam ii1082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1083 ( .DX(\a_dinx[6]_cal1_u146_mac ), .F0(\c1r1_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1083.CONFIG_DATA = 16'hCA00;
      defparam ii1083.PLACE_LOCATION = "NONE";
      defparam ii1083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1084 ( .DX(\a_dinx[6]_cal1_u147_mac ), .F0(\c1r1_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1084.CONFIG_DATA = 16'hCA00;
      defparam ii1084.PLACE_LOCATION = "NONE";
      defparam ii1084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1085 ( .DX(nn1085), .F0(\c1r1_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_149_) );
      defparam ii1085.CONFIG_DATA = 16'hCACA;
      defparam ii1085.PLACE_LOCATION = "NONE";
      defparam ii1085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1086 ( .DX(\a_dinx[6]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u146_mac ), .F3(nn1085) );
      defparam ii1086.CONFIG_DATA = 16'hE4A0;
      defparam ii1086.PLACE_LOCATION = "NONE";
      defparam ii1086.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1087 ( .DX(nn1087), .F0(\c1r1_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r3_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_150_) );
      defparam ii1087.CONFIG_DATA = 16'hCACA;
      defparam ii1087.PLACE_LOCATION = "NONE";
      defparam ii1087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1088 ( .DX(\a_dinx[6]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[6]_cal1_u147_mac ), .F3(nn1087) );
      defparam ii1088.CONFIG_DATA = 16'hE4A0;
      defparam ii1088.PLACE_LOCATION = "NONE";
      defparam ii1088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1089 ( .DX(\a_dinx[7]_cal1_u138_mac ), .F0(\c1r1_q[3]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1089.CONFIG_DATA = 16'hCA00;
      defparam ii1089.PLACE_LOCATION = "NONE";
      defparam ii1089.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1090 ( .DX(\a_dinx[7]_cal1_u139_mac ), .F0(\c1r1_q[12]_fifo1_ram_inst_0A_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_0A_u_emb18k_1 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1090.CONFIG_DATA = 16'hCA00;
      defparam ii1090.PLACE_LOCATION = "NONE";
      defparam ii1090.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1091 ( .DX(nn1091), .F0(\c1r1_q[3]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[3]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_151_) );
      defparam ii1091.CONFIG_DATA = 16'hCACA;
      defparam ii1091.PLACE_LOCATION = "NONE";
      defparam ii1091.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1092 ( .DX(\a_dinx[7]_cal1_u140_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u138_mac ), .F3(nn1091) );
      defparam ii1092.CONFIG_DATA = 16'hE4A0;
      defparam ii1092.PLACE_LOCATION = "NONE";
      defparam ii1092.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1093 ( .DX(nn1093), .F0(\c1r1_q[12]_fifo1_ram_inst_1A_u_emb18k_1 ), .F1(\c1r3_q[12]_fifo1_ram_inst_1A_u_emb18k_1 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_152_) );
      defparam ii1093.CONFIG_DATA = 16'hCACA;
      defparam ii1093.PLACE_LOCATION = "NONE";
      defparam ii1093.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1094 ( .DX(\a_dinx[7]_cal1_u141_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u139_mac ), .F3(nn1093) );
      defparam ii1094.CONFIG_DATA = 16'hE4A0;
      defparam ii1094.PLACE_LOCATION = "NONE";
      defparam ii1094.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1095 ( .DX(\a_dinx[7]_cal1_u142_mac ), .F0(\c1r1_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1095.CONFIG_DATA = 16'hCA00;
      defparam ii1095.PLACE_LOCATION = "NONE";
      defparam ii1095.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1096 ( .DX(\a_dinx[7]_cal1_u143_mac ), .F0(\c1r1_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_0A_u_emb18k_0 ), .F2(\fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1096.CONFIG_DATA = 16'hCA00;
      defparam ii1096.PLACE_LOCATION = "NONE";
      defparam ii1096.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1097 ( .DX(nn1097), .F0(\c1r1_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[1]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_153_) );
      defparam ii1097.CONFIG_DATA = 16'hCACA;
      defparam ii1097.PLACE_LOCATION = "NONE";
      defparam ii1097.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1098 ( .DX(\a_dinx[7]_cal1_u144_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u142_mac ), .F3(nn1097) );
      defparam ii1098.CONFIG_DATA = 16'hE4A0;
      defparam ii1098.PLACE_LOCATION = "NONE";
      defparam ii1098.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1099 ( .DX(nn1099), .F0(\c1r1_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ), .F1(\c1r3_q[10]_fifo1_ram_inst_1A_u_emb18k_0 ), .F2(\fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_154_) );
      defparam ii1099.CONFIG_DATA = 16'hCACA;
      defparam ii1099.PLACE_LOCATION = "NONE";
      defparam ii1099.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1100 ( .DX(\a_dinx[7]_cal1_u145_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u143_mac ), .F3(nn1099) );
      defparam ii1100.CONFIG_DATA = 16'hE4A0;
      defparam ii1100.PLACE_LOCATION = "NONE";
      defparam ii1100.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1101 ( .DX(\a_dinx[7]_cal1_u146_mac ), .F0(\c1r2_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1101.CONFIG_DATA = 16'hCA00;
      defparam ii1101.PLACE_LOCATION = "NONE";
      defparam ii1101.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1102 ( .DX(\a_dinx[7]_cal1_u147_mac ), .F0(\c1r2_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_0B_u_emb18k_0 ), .F2(\fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net ), .F3(nn0882) );
      defparam ii1102.CONFIG_DATA = 16'hCA00;
      defparam ii1102.PLACE_LOCATION = "NONE";
      defparam ii1102.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1103 ( .DX(nn1103), .F0(\c1r2_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[2]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net ), .F3(dummy_abc_155_) );
      defparam ii1103.CONFIG_DATA = 16'hCACA;
      defparam ii1103.PLACE_LOCATION = "NONE";
      defparam ii1103.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1104 ( .DX(\a_dinx[7]_cal1_u148_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u146_mac ), .F3(nn1103) );
      defparam ii1104.CONFIG_DATA = 16'hE4A0;
      defparam ii1104.PLACE_LOCATION = "NONE";
      defparam ii1104.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1105 ( .DX(nn1105), .F0(\c1r2_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ), .F1(\c1r4_q[11]_fifo1_ram_inst_1B_u_emb18k_0 ), .F2(\fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net ), .F3(dummy_abc_156_) );
      defparam ii1105.CONFIG_DATA = 16'hCACA;
      defparam ii1105.PLACE_LOCATION = "NONE";
      defparam ii1105.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1106 ( .DX(\a_dinx[7]_cal1_u149_mac ), .F0(dummy_62_), .F1(nn0882), .F2(\a_dinx[7]_cal1_u147_mac ), .F3(nn1105) );
      defparam ii1106.CONFIG_DATA = 16'hE4A0;
      defparam ii1106.PLACE_LOCATION = "NONE";
      defparam ii1106.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1107 ( .DX(nn1107), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[0]|Q_net ), .F2(\cal1_v__reg[0]|Q_net ), .F3(dummy_abc_157_) );
      defparam ii1107.CONFIG_DATA = 16'h9696;
      defparam ii1107.PLACE_LOCATION = "NONE";
      defparam ii1107.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1108 ( .DX(nn1108), .F0(\cal1_uPreF__reg[0]|Q_net ), .F1(dummy_abc_158_), .F2(dummy_abc_159_), .F3(dummy_abc_160_) );
      defparam ii1108.CONFIG_DATA = 16'h5555;
      defparam ii1108.PLACE_LOCATION = "NONE";
      defparam ii1108.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1109 ( .DX(nn1109), .F0(\cal1_uPreF__reg[1]|Q_net ), .F1(dummy_abc_161_), .F2(dummy_abc_162_), .F3(dummy_abc_163_) );
      defparam ii1109.CONFIG_DATA = 16'h5555;
      defparam ii1109.PLACE_LOCATION = "NONE";
      defparam ii1109.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1110 ( .DX(nn1110), .F0(\cal1_uPreF__reg[2]|Q_net ), .F1(dummy_abc_164_), .F2(dummy_abc_165_), .F3(dummy_abc_166_) );
      defparam ii1110.CONFIG_DATA = 16'h5555;
      defparam ii1110.PLACE_LOCATION = "NONE";
      defparam ii1110.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1111 ( .DX(nn1111), .F0(\cal1_uPreF__reg[3]|Q_net ), .F1(dummy_abc_167_), .F2(dummy_abc_168_), .F3(dummy_abc_169_) );
      defparam ii1111.CONFIG_DATA = 16'h5555;
      defparam ii1111.PLACE_LOCATION = "NONE";
      defparam ii1111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1112 ( .DX(nn1112), .F0(\cal1_uPreF__reg[4]|Q_net ), .F1(dummy_abc_170_), .F2(dummy_abc_171_), .F3(dummy_abc_172_) );
      defparam ii1112.CONFIG_DATA = 16'h5555;
      defparam ii1112.PLACE_LOCATION = "NONE";
      defparam ii1112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1113 ( .DX(nn1113), .F0(\cal1_uPreF__reg[5]|Q_net ), .F1(dummy_abc_173_), .F2(dummy_abc_174_), .F3(dummy_abc_175_) );
      defparam ii1113.CONFIG_DATA = 16'h5555;
      defparam ii1113.PLACE_LOCATION = "NONE";
      defparam ii1113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1114 ( .DX(nn1114), .F0(dummy_abc_176_), .F1(dummy_abc_177_), .F2(dummy_abc_178_), .F3(dummy_abc_179_) );
      defparam ii1114.CONFIG_DATA = 16'h0000;
      defparam ii1114.PLACE_LOCATION = "NONE";
      defparam ii1114.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7_209_ ( 
        .CA( {a_dinxy_cen_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_885_ ), 
        .DX( {nn1114, nn1113, nn1112, nn1111, nn1110, nn1109, nn1108} ), 
        .SUM( {\cal1_u54_XORCI_6|SUM_net , \cal1_u54_XORCI_5|SUM_net , 
              \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_3|SUM_net , \cal1_u54_XORCI_2|SUM_net , 
              \cal1_u54_XORCI_1|SUM_net , \cal1_u54_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1124 ( .DX(nn1124), .F0(\cal1_uPreF__reg[0]|Q_net ), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_abc_180_), .F3(dummy_abc_181_) );
      defparam ii1124.CONFIG_DATA = 16'h9999;
      defparam ii1124.PLACE_LOCATION = "NONE";
      defparam ii1124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1125 ( .DX(nn1125), .F0(\cal1_v__reg[1]|Q_net ), .F1(\cal1_u54_XORCI_1|SUM_net ), .F2(dummy_abc_182_), .F3(dummy_abc_183_) );
      defparam ii1125.CONFIG_DATA = 16'h9999;
      defparam ii1125.PLACE_LOCATION = "NONE";
      defparam ii1125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1126 ( .DX(nn1126), .F0(\cal1_v__reg[2]|Q_net ), .F1(\cal1_u54_XORCI_2|SUM_net ), .F2(dummy_abc_184_), .F3(dummy_abc_185_) );
      defparam ii1126.CONFIG_DATA = 16'h9999;
      defparam ii1126.PLACE_LOCATION = "NONE";
      defparam ii1126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1127 ( .DX(nn1127), .F0(\cal1_v__reg[3]|Q_net ), .F1(\cal1_u54_XORCI_3|SUM_net ), .F2(dummy_abc_186_), .F3(dummy_abc_187_) );
      defparam ii1127.CONFIG_DATA = 16'h9999;
      defparam ii1127.PLACE_LOCATION = "NONE";
      defparam ii1127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1128 ( .DX(nn1128), .F0(\cal1_v__reg[4]|Q_net ), .F1(\cal1_u54_XORCI_4|SUM_net ), .F2(dummy_abc_188_), .F3(dummy_abc_189_) );
      defparam ii1128.CONFIG_DATA = 16'h9999;
      defparam ii1128.PLACE_LOCATION = "NONE";
      defparam ii1128.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1129 ( .DX(nn1129), .F0(\cal1_v__reg[5]|Q_net ), .F1(\cal1_u54_XORCI_5|SUM_net ), .F2(dummy_abc_190_), .F3(dummy_abc_191_) );
      defparam ii1129.CONFIG_DATA = 16'h9999;
      defparam ii1129.PLACE_LOCATION = "NONE";
      defparam ii1129.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1130 ( .DX(nn1130), .F0(\cal1_u54_XORCI_6|SUM_net ), .F1(dummy_abc_192_), .F2(dummy_abc_193_), .F3(dummy_abc_194_) );
      defparam ii1130.CONFIG_DATA = 16'h5555;
      defparam ii1130.PLACE_LOCATION = "NONE";
      defparam ii1130.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7_210_ ( 
        .CA( {\cal1_u54_XORCI_6|SUM_net , \cal1_u54_XORCI_5|SUM_net , 
              \cal1_u54_XORCI_4|SUM_net , \cal1_u54_XORCI_3|SUM_net , \cal1_u54_XORCI_2|SUM_net , 
              \cal1_u54_XORCI_1|SUM_net , \cal1_uPreF__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_886_ ), 
        .DX( {nn1130, nn1129, nn1128, nn1127, nn1126, nn1125, nn1124} ), 
        .SUM( {\cal1_u55_XORCI_6|SUM_net , \cal1_u55_XORCI_5|SUM_net , 
              \cal1_u55_XORCI_4|SUM_net , \cal1_u55_XORCI_3|SUM_net , \cal1_u55_XORCI_2|SUM_net , 
              \cal1_u55_XORCI_1|SUM_net , \cal1_u55_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1140 ( .DX(nn1140), .F0(\a_mac_out[7]_cal1_u137_mac ), .F1(\cal1_u55_XORCI_1|SUM_net ), .F2(dummy_abc_195_), .F3(dummy_abc_196_) );
      defparam ii1140.CONFIG_DATA = 16'h6666;
      defparam ii1140.PLACE_LOCATION = "NONE";
      defparam ii1140.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1141 ( .DX(nn1141), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\cal1_u55_XORCI_2|SUM_net ), .F2(dummy_abc_197_), .F3(dummy_abc_198_) );
      defparam ii1141.CONFIG_DATA = 16'h6666;
      defparam ii1141.PLACE_LOCATION = "NONE";
      defparam ii1141.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1142 ( .DX(nn1142), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(\cal1_u55_XORCI_3|SUM_net ), .F2(dummy_abc_199_), .F3(dummy_abc_200_) );
      defparam ii1142.CONFIG_DATA = 16'h6666;
      defparam ii1142.PLACE_LOCATION = "NONE";
      defparam ii1142.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1143 ( .DX(nn1143), .F0(\a_mac_out[10]_cal1_u137_mac ), .F1(\cal1_u55_XORCI_4|SUM_net ), .F2(dummy_abc_201_), .F3(dummy_abc_202_) );
      defparam ii1143.CONFIG_DATA = 16'h6666;
      defparam ii1143.PLACE_LOCATION = "NONE";
      defparam ii1143.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1144 ( .DX(nn1144), .F0(\a_mac_out[11]_cal1_u137_mac ), .F1(\cal1_u55_XORCI_5|SUM_net ), .F2(dummy_abc_203_), .F3(dummy_abc_204_) );
      defparam ii1144.CONFIG_DATA = 16'h6666;
      defparam ii1144.PLACE_LOCATION = "NONE";
      defparam ii1144.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1145 ( .DX(nn1145), .F0(\cal1_u55_XORCI_6|SUM_net ), .F1(dummy_abc_205_), .F2(dummy_abc_206_), .F3(dummy_abc_207_) );
      defparam ii1145.CONFIG_DATA = 16'hAAAA;
      defparam ii1145.PLACE_LOCATION = "NONE";
      defparam ii1145.PCK_LOCATION = "NONE";
    scaler_ipc_adder_7 carry_7 ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[11]_cal1_u137_mac , 
              \a_mac_out[10]_cal1_u137_mac , \a_mac_out[9]_cal1_u137_mac , \a_mac_out[8]_cal1_u137_mac , 
              \a_mac_out[7]_cal1_u137_mac , \a_mac_out[6]_cal1_u137_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_884_ ), 
        .DX( {nn1145, nn1144, nn1143, nn1142, nn1141, nn1140, nn1107} ), 
        .SUM( {\cal1_u133_XORCI_6|SUM_net , \cal1_u133_XORCI_5|SUM_net , 
              \cal1_u133_XORCI_4|SUM_net , \cal1_u133_XORCI_3|SUM_net , \cal1_u133_XORCI_2|SUM_net , 
              \cal1_u133_XORCI_1|SUM_net , \cal1_u133_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1155 ( .DX(\a_diny[0]_cal1_u139_mac ), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[0]|Q_net ), .F2(dummy_abc_208_), .F3(dummy_abc_209_) );
      defparam ii1155.CONFIG_DATA = 16'h6666;
      defparam ii1155.PLACE_LOCATION = "NONE";
      defparam ii1155.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1156 ( .DX(\a_diny[0]_cal1_u140_mac ), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\cal1_v__reg[0]|Q_net ), .F2(dummy_abc_210_), .F3(dummy_abc_211_) );
      defparam ii1156.CONFIG_DATA = 16'h6666;
      defparam ii1156.PLACE_LOCATION = "NONE";
      defparam ii1156.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1157 ( .DX(\a_diny[1]_cal1_u139_mac ), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\a_mac_out[7]_cal1_u137_mac ), .F2(\cal1_uPreF__reg[0]|Q_net ), .F3(\cal1_uPreF__reg[1]|Q_net ) );
      defparam ii1157.CONFIG_DATA = 16'h39C6;
      defparam ii1157.PLACE_LOCATION = "NONE";
      defparam ii1157.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1158 ( .DX(\a_diny[1]_cal1_u140_mac ), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\a_mac_out[7]_cal1_u137_mac ), .F2(\cal1_v__reg[0]|Q_net ), .F3(\cal1_v__reg[1]|Q_net ) );
      defparam ii1158.CONFIG_DATA = 16'h39C6;
      defparam ii1158.PLACE_LOCATION = "NONE";
      defparam ii1158.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1159 ( .DX(nn1159), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\a_mac_out[7]_cal1_u137_mac ), .F2(\cal1_uPreF__reg[0]|Q_net ), .F3(\cal1_uPreF__reg[1]|Q_net ) );
      defparam ii1159.CONFIG_DATA = 16'hF731;
      defparam ii1159.PLACE_LOCATION = "NONE";
      defparam ii1159.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1160 ( .DX(\a_diny[2]_cal1_u139_mac ), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[2]|Q_net ), .F2(nn1159), .F3(dummy_abc_212_) );
      defparam ii1160.CONFIG_DATA = 16'h6969;
      defparam ii1160.PLACE_LOCATION = "NONE";
      defparam ii1160.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1161 ( .DX(nn1161), .F0(\a_mac_out[6]_cal1_u137_mac ), .F1(\a_mac_out[7]_cal1_u137_mac ), .F2(\cal1_v__reg[0]|Q_net ), .F3(\cal1_v__reg[1]|Q_net ) );
      defparam ii1161.CONFIG_DATA = 16'hF731;
      defparam ii1161.PLACE_LOCATION = "NONE";
      defparam ii1161.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1162 ( .DX(\a_diny[2]_cal1_u140_mac ), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\cal1_v__reg[2]|Q_net ), .F2(nn1161), .F3(dummy_abc_213_) );
      defparam ii1162.CONFIG_DATA = 16'h6969;
      defparam ii1162.PLACE_LOCATION = "NONE";
      defparam ii1162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1163 ( .DX(nn1163), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[2]|Q_net ), .F2(nn1159), .F3(dummy_abc_214_) );
      defparam ii1163.CONFIG_DATA = 16'h2B2B;
      defparam ii1163.PLACE_LOCATION = "NONE";
      defparam ii1163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1164 ( .DX(\a_diny[3]_cal1_u139_mac ), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[3]|Q_net ), .F2(nn1163), .F3(dummy_abc_215_) );
      defparam ii1164.CONFIG_DATA = 16'h9696;
      defparam ii1164.PLACE_LOCATION = "NONE";
      defparam ii1164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1165 ( .DX(nn1165), .F0(\a_mac_out[8]_cal1_u137_mac ), .F1(\cal1_v__reg[2]|Q_net ), .F2(nn1161), .F3(dummy_abc_216_) );
      defparam ii1165.CONFIG_DATA = 16'h2B2B;
      defparam ii1165.PLACE_LOCATION = "NONE";
      defparam ii1165.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1166 ( .DX(\a_diny[3]_cal1_u140_mac ), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(\cal1_v__reg[3]|Q_net ), .F2(nn1165), .F3(dummy_abc_217_) );
      defparam ii1166.CONFIG_DATA = 16'h9696;
      defparam ii1166.PLACE_LOCATION = "NONE";
      defparam ii1166.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1167 ( .DX(nn1167), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[3]|Q_net ), .F2(nn1163), .F3(dummy_abc_218_) );
      defparam ii1167.CONFIG_DATA = 16'h4D4D;
      defparam ii1167.PLACE_LOCATION = "NONE";
      defparam ii1167.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1168 ( .DX(\a_diny[4]_cal1_u139_mac ), .F0(\a_mac_out[10]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[4]|Q_net ), .F2(nn1167), .F3(dummy_abc_219_) );
      defparam ii1168.CONFIG_DATA = 16'h6969;
      defparam ii1168.PLACE_LOCATION = "NONE";
      defparam ii1168.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1169 ( .DX(nn1169), .F0(\a_mac_out[9]_cal1_u137_mac ), .F1(\cal1_v__reg[3]|Q_net ), .F2(nn1165), .F3(dummy_abc_220_) );
      defparam ii1169.CONFIG_DATA = 16'h4D4D;
      defparam ii1169.PLACE_LOCATION = "NONE";
      defparam ii1169.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1170 ( .DX(\a_diny[4]_cal1_u140_mac ), .F0(\a_mac_out[10]_cal1_u137_mac ), .F1(\cal1_v__reg[4]|Q_net ), .F2(nn1169), .F3(dummy_abc_221_) );
      defparam ii1170.CONFIG_DATA = 16'h6969;
      defparam ii1170.PLACE_LOCATION = "NONE";
      defparam ii1170.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1171 ( .DX(nn1171), .F0(\a_mac_out[11]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[5]|Q_net ), .F2(dummy_abc_222_), .F3(dummy_abc_223_) );
      defparam ii1171.CONFIG_DATA = 16'h6666;
      defparam ii1171.PLACE_LOCATION = "NONE";
      defparam ii1171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1172 ( .DX(\a_diny[5]_cal1_u139_mac ), .F0(\a_mac_out[10]_cal1_u137_mac ), .F1(\cal1_uPreF__reg[4]|Q_net ), .F2(nn1167), .F3(nn1171) );
      defparam ii1172.CONFIG_DATA = 16'hD42B;
      defparam ii1172.PLACE_LOCATION = "NONE";
      defparam ii1172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1173 ( .DX(nn1173), .F0(\a_mac_out[11]_cal1_u137_mac ), .F1(\cal1_v__reg[5]|Q_net ), .F2(dummy_abc_224_), .F3(dummy_abc_225_) );
      defparam ii1173.CONFIG_DATA = 16'h6666;
      defparam ii1173.PLACE_LOCATION = "NONE";
      defparam ii1173.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1174 ( .DX(\a_diny[5]_cal1_u140_mac ), .F0(\a_mac_out[10]_cal1_u137_mac ), .F1(\cal1_v__reg[4]|Q_net ), .F2(nn1169), .F3(nn1173) );
      defparam ii1174.CONFIG_DATA = 16'hD42B;
      defparam ii1174.PLACE_LOCATION = "NONE";
      defparam ii1174.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1175 ( .DX(u8231_O), .F0(rst), .F1(u5859_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(dummy_abc_226_) );
      defparam ii1175.CONFIG_DATA = 16'hEAEA;
      defparam ii1175.PLACE_LOCATION = "NONE";
      defparam ii1175.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1176 ( .DX(\c1r1_aa[10]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F2(u8231_O), .F3(dummy_abc_227_) );
      defparam ii1176.CONFIG_DATA = 16'hCACA;
      defparam ii1176.PLACE_LOCATION = "NONE";
      defparam ii1176.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1177 ( .DX(\c1r1_aa[10]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[8]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F3(u8231_O) );
      defparam ii1177.CONFIG_DATA = 16'hD8CC;
      defparam ii1177.PLACE_LOCATION = "NONE";
      defparam ii1177.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1178 ( .DX(\c1r1_aa[11]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F2(u8231_O), .F3(dummy_abc_228_) );
      defparam ii1178.CONFIG_DATA = 16'hCACA;
      defparam ii1178.PLACE_LOCATION = "NONE";
      defparam ii1178.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1179 ( .DX(\c1r1_aa[11]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[9]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F3(u8231_O) );
      defparam ii1179.CONFIG_DATA = 16'hD8CC;
      defparam ii1179.PLACE_LOCATION = "NONE";
      defparam ii1179.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1180 ( .DX(\c1r1_aa[2]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F2(u8231_O), .F3(dummy_abc_229_) );
      defparam ii1180.CONFIG_DATA = 16'hCACA;
      defparam ii1180.PLACE_LOCATION = "NONE";
      defparam ii1180.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1181 ( .DX(\c1r1_aa[2]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[0]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F3(u8231_O) );
      defparam ii1181.CONFIG_DATA = 16'hD8CC;
      defparam ii1181.PLACE_LOCATION = "NONE";
      defparam ii1181.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1182 ( .DX(\c1r1_aa[3]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F2(u8231_O), .F3(dummy_abc_230_) );
      defparam ii1182.CONFIG_DATA = 16'hCACA;
      defparam ii1182.PLACE_LOCATION = "NONE";
      defparam ii1182.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1183 ( .DX(\c1r1_aa[3]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[1]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F3(u8231_O) );
      defparam ii1183.CONFIG_DATA = 16'hD8CC;
      defparam ii1183.PLACE_LOCATION = "NONE";
      defparam ii1183.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1184 ( .DX(\c1r1_aa[4]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F2(u8231_O), .F3(dummy_abc_231_) );
      defparam ii1184.CONFIG_DATA = 16'hCACA;
      defparam ii1184.PLACE_LOCATION = "NONE";
      defparam ii1184.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1185 ( .DX(\c1r1_aa[4]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[2]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F3(u8231_O) );
      defparam ii1185.CONFIG_DATA = 16'hD8CC;
      defparam ii1185.PLACE_LOCATION = "NONE";
      defparam ii1185.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1186 ( .DX(\c1r1_aa[5]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F2(u8231_O), .F3(dummy_abc_232_) );
      defparam ii1186.CONFIG_DATA = 16'hCACA;
      defparam ii1186.PLACE_LOCATION = "NONE";
      defparam ii1186.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1187 ( .DX(\c1r1_aa[5]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[3]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F3(u8231_O) );
      defparam ii1187.CONFIG_DATA = 16'hD8CC;
      defparam ii1187.PLACE_LOCATION = "NONE";
      defparam ii1187.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1188 ( .DX(\c1r1_aa[6]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F2(u8231_O), .F3(dummy_abc_233_) );
      defparam ii1188.CONFIG_DATA = 16'hCACA;
      defparam ii1188.PLACE_LOCATION = "NONE";
      defparam ii1188.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1189 ( .DX(\c1r1_aa[6]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[4]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F3(u8231_O) );
      defparam ii1189.CONFIG_DATA = 16'hD8CC;
      defparam ii1189.PLACE_LOCATION = "NONE";
      defparam ii1189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1190 ( .DX(\c1r1_aa[7]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F2(u8231_O), .F3(dummy_abc_234_) );
      defparam ii1190.CONFIG_DATA = 16'hCACA;
      defparam ii1190.PLACE_LOCATION = "NONE";
      defparam ii1190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1191 ( .DX(\c1r1_aa[7]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[5]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F3(u8231_O) );
      defparam ii1191.CONFIG_DATA = 16'hD8CC;
      defparam ii1191.PLACE_LOCATION = "NONE";
      defparam ii1191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1192 ( .DX(\c1r1_aa[8]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F2(u8231_O), .F3(dummy_abc_235_) );
      defparam ii1192.CONFIG_DATA = 16'hCACA;
      defparam ii1192.PLACE_LOCATION = "NONE";
      defparam ii1192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1193 ( .DX(\c1r1_aa[8]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[6]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F3(u8231_O) );
      defparam ii1193.CONFIG_DATA = 16'hD8CC;
      defparam ii1193.PLACE_LOCATION = "NONE";
      defparam ii1193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1194 ( .DX(\c1r1_aa[9]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F2(u8231_O), .F3(dummy_abc_236_) );
      defparam ii1194.CONFIG_DATA = 16'hCACA;
      defparam ii1194.PLACE_LOCATION = "NONE";
      defparam ii1194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1195 ( .DX(\c1r1_aa[9]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[7]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F3(u8231_O) );
      defparam ii1195.CONFIG_DATA = 16'hD8CC;
      defparam ii1195.PLACE_LOCATION = "NONE";
      defparam ii1195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1196 ( .DX(nn1196), .F0(\cal1_u__reg[11]|Q_net ), .F1(nn0886), .F2(dummy_abc_237_), .F3(dummy_abc_238_) );
      defparam ii1196.CONFIG_DATA = 16'h6666;
      defparam ii1196.PLACE_LOCATION = "NONE";
      defparam ii1196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1197 ( .DX(nn1197), .F0(\cal1_u__reg[12]|Q_net ), .F1(\u3_XORCI_1|SUM_net ), .F2(dummy_abc_239_), .F3(dummy_abc_240_) );
      defparam ii1197.CONFIG_DATA = 16'h9999;
      defparam ii1197.PLACE_LOCATION = "NONE";
      defparam ii1197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1198 ( .DX(nn1198), .F0(\cal1_u__reg[13]|Q_net ), .F1(\u3_XORCI_2|SUM_net ), .F2(dummy_abc_241_), .F3(dummy_abc_242_) );
      defparam ii1198.CONFIG_DATA = 16'h9999;
      defparam ii1198.PLACE_LOCATION = "NONE";
      defparam ii1198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1199 ( .DX(nn1199), .F0(\cal1_u__reg[14]|Q_net ), .F1(\u3_XORCI_3|SUM_net ), .F2(dummy_abc_243_), .F3(dummy_abc_244_) );
      defparam ii1199.CONFIG_DATA = 16'h9999;
      defparam ii1199.PLACE_LOCATION = "NONE";
      defparam ii1199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1200 ( .DX(nn1200), .F0(\cal1_u__reg[15]|Q_net ), .F1(\u3_XORCI_4|SUM_net ), .F2(dummy_abc_245_), .F3(dummy_abc_246_) );
      defparam ii1200.CONFIG_DATA = 16'h9999;
      defparam ii1200.PLACE_LOCATION = "NONE";
      defparam ii1200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1201 ( .DX(nn1201), .F0(\cal1_u__reg[16]|Q_net ), .F1(\u3_XORCI_5|SUM_net ), .F2(dummy_abc_247_), .F3(dummy_abc_248_) );
      defparam ii1201.CONFIG_DATA = 16'h9999;
      defparam ii1201.PLACE_LOCATION = "NONE";
      defparam ii1201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1202 ( .DX(nn1202), .F0(\u3_XORCI_6|SUM_net ), .F1(dummy_abc_249_), .F2(dummy_abc_250_), .F3(dummy_abc_251_) );
      defparam ii1202.CONFIG_DATA = 16'h5555;
      defparam ii1202.PLACE_LOCATION = "NONE";
      defparam ii1202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1203 ( .DX(nn1203), .F0(\u3_XORCI_7|SUM_net ), .F1(dummy_abc_252_), .F2(dummy_abc_253_), .F3(dummy_abc_254_) );
      defparam ii1203.CONFIG_DATA = 16'h5555;
      defparam ii1203.PLACE_LOCATION = "NONE";
      defparam ii1203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1204 ( .DX(nn1204), .F0(\u3_XORCI_8|SUM_net ), .F1(dummy_abc_255_), .F2(dummy_abc_256_), .F3(dummy_abc_257_) );
      defparam ii1204.CONFIG_DATA = 16'h5555;
      defparam ii1204.PLACE_LOCATION = "NONE";
      defparam ii1204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1205 ( .DX(nn1205), .F0(\u3_XORCI_9|SUM_net ), .F1(dummy_abc_258_), .F2(dummy_abc_259_), .F3(dummy_abc_260_) );
      defparam ii1205.CONFIG_DATA = 16'h5555;
      defparam ii1205.PLACE_LOCATION = "NONE";
      defparam ii1205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1206 ( .DX(nn1206), .F0(\u3_XORCI_10|SUM_net ), .F1(dummy_abc_261_), .F2(dummy_abc_262_), .F3(dummy_abc_263_) );
      defparam ii1206.CONFIG_DATA = 16'h5555;
      defparam ii1206.PLACE_LOCATION = "NONE";
      defparam ii1206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1207 ( .DX(nn1207), .F0(dummy_abc_264_), .F1(dummy_abc_265_), .F2(dummy_abc_266_), .F3(dummy_abc_267_) );
      defparam ii1207.CONFIG_DATA = 16'hFFFF;
      defparam ii1207.PLACE_LOCATION = "NONE";
      defparam ii1207.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_212_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, \cal1_u__reg[16]|Q_net , \cal1_u__reg[15]|Q_net , 
              \cal1_u__reg[14]|Q_net , \cal1_u__reg[13]|Q_net , \cal1_u__reg[12]|Q_net , 
              \cal1_u__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_49_ ), 
        .DX( {nn1207, nn1206, nn1205, nn1204, nn1203, nn1202, nn1201, nn1200, 
              nn1199, nn1198, nn1197, nn1196} ), 
        .SUM( {\cal1_u61_XORCI_11|SUM_net , dummy_50_, dummy_51_, dummy_52_, 
              dummy_53_, dummy_54_, dummy_55_, dummy_56_, dummy_57_, dummy_58_, 
              dummy_59_, dummy_60_} )
      );
    CS_LUT4_PRIM ii1222 ( .DX(nn1222), .F0(dummy_49_), .F1(dummy_abc_268_), .F2(dummy_abc_269_), .F3(dummy_abc_270_) );
      defparam ii1222.CONFIG_DATA = 16'h5555;
      defparam ii1222.PLACE_LOCATION = "NONE";
      defparam ii1222.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1223 ( .DX(nn1223), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(dummy_49_), .F2(dummy_abc_271_), .F3(dummy_abc_272_) );
      defparam ii1223.CONFIG_DATA = 16'h9999;
      defparam ii1223.PLACE_LOCATION = "NONE";
      defparam ii1223.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1224 ( .DX(nn1224), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(dummy_abc_273_), .F2(dummy_abc_274_), .F3(dummy_abc_275_) );
      defparam ii1224.CONFIG_DATA = 16'hAAAA;
      defparam ii1224.PLACE_LOCATION = "NONE";
      defparam ii1224.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1225 ( .DX(nn1225), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(dummy_abc_276_), .F2(dummy_abc_277_), .F3(dummy_abc_278_) );
      defparam ii1225.CONFIG_DATA = 16'hAAAA;
      defparam ii1225.PLACE_LOCATION = "NONE";
      defparam ii1225.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1226 ( .DX(nn1226), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(dummy_abc_279_), .F2(dummy_abc_280_), .F3(dummy_abc_281_) );
      defparam ii1226.CONFIG_DATA = 16'hAAAA;
      defparam ii1226.PLACE_LOCATION = "NONE";
      defparam ii1226.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1227 ( .DX(nn1227), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(dummy_abc_282_), .F2(dummy_abc_283_), .F3(dummy_abc_284_) );
      defparam ii1227.CONFIG_DATA = 16'hAAAA;
      defparam ii1227.PLACE_LOCATION = "NONE";
      defparam ii1227.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1228 ( .DX(nn1228), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(dummy_abc_285_), .F2(dummy_abc_286_), .F3(dummy_abc_287_) );
      defparam ii1228.CONFIG_DATA = 16'hAAAA;
      defparam ii1228.PLACE_LOCATION = "NONE";
      defparam ii1228.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1229 ( .DX(nn1229), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(dummy_abc_288_), .F2(dummy_abc_289_), .F3(dummy_abc_290_) );
      defparam ii1229.CONFIG_DATA = 16'hAAAA;
      defparam ii1229.PLACE_LOCATION = "NONE";
      defparam ii1229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1230 ( .DX(nn1230), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(dummy_abc_291_), .F2(dummy_abc_292_), .F3(dummy_abc_293_) );
      defparam ii1230.CONFIG_DATA = 16'hAAAA;
      defparam ii1230.PLACE_LOCATION = "NONE";
      defparam ii1230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1231 ( .DX(nn1231), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(dummy_abc_294_), .F2(dummy_abc_295_), .F3(dummy_abc_296_) );
      defparam ii1231.CONFIG_DATA = 16'hAAAA;
      defparam ii1231.PLACE_LOCATION = "NONE";
      defparam ii1231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1232 ( .DX(nn1232), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(dummy_abc_297_), .F2(dummy_abc_298_), .F3(dummy_abc_299_) );
      defparam ii1232.CONFIG_DATA = 16'hAAAA;
      defparam ii1232.PLACE_LOCATION = "NONE";
      defparam ii1232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1233 ( .DX(nn1233), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(dummy_abc_300_), .F2(dummy_abc_301_), .F3(dummy_abc_302_) );
      defparam ii1233.CONFIG_DATA = 16'hAAAA;
      defparam ii1233.PLACE_LOCATION = "NONE";
      defparam ii1233.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11 ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn1222} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_13_ ), 
        .DX( {nn1233, nn1232, nn1231, nn1230, nn1229, nn1228, nn1227, nn1226, 
              nn1225, nn1224, nn1223} ), 
        .SUM( {\cal1_u129_XORCI_10|SUM_net , \cal1_u129_XORCI_9|SUM_net , 
              \cal1_u129_XORCI_8|SUM_net , \cal1_u129_XORCI_7|SUM_net , \cal1_u129_XORCI_6|SUM_net , 
              \cal1_u129_XORCI_5|SUM_net , \cal1_u129_XORCI_4|SUM_net , \cal1_u129_XORCI_3|SUM_net , 
              \cal1_u129_XORCI_2|SUM_net , \cal1_u129_XORCI_1|SUM_net , \cal1_u129_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1247 ( .DX(c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0), .F0(clka), .F1(clkb), .F2(u8231_O), .F3(dummy_abc_303_) );
      defparam ii1247.CONFIG_DATA = 16'hACAC;
      defparam ii1247.PLACE_LOCATION = "NONE";
      defparam ii1247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1248 ( .DX(c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0), .F0(clka), .F1(clkb), .F2(rst), .F3(u8231_O) );
      defparam ii1248.CONFIG_DATA = 16'hCACC;
      defparam ii1248.PLACE_LOCATION = "NONE";
      defparam ii1248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1249 ( .DX(nn1249), .F0(\a_mac_out[6]_cal1_u148_mac ), .F1(\a_mac_out[6]_cal1_u149_mac ), .F2(dummy_abc_304_), .F3(dummy_abc_305_) );
      defparam ii1249.CONFIG_DATA = 16'h6666;
      defparam ii1249.PLACE_LOCATION = "NONE";
      defparam ii1249.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1250 ( .DX(nn1250), .F0(\a_mac_out[6]_cal1_u148_mac ), .F1(\a_mac_out[6]_cal1_u149_mac ), .F2(dummy_abc_306_), .F3(dummy_abc_307_) );
      defparam ii1250.CONFIG_DATA = 16'h6666;
      defparam ii1250.PLACE_LOCATION = "NONE";
      defparam ii1250.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1251 ( .DX(nn1251), .F0(\a_mac_out[7]_cal1_u148_mac ), .F1(\a_mac_out[7]_cal1_u149_mac ), .F2(dummy_abc_308_), .F3(dummy_abc_309_) );
      defparam ii1251.CONFIG_DATA = 16'h6666;
      defparam ii1251.PLACE_LOCATION = "NONE";
      defparam ii1251.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1252 ( .DX(nn1252), .F0(\a_mac_out[8]_cal1_u148_mac ), .F1(\a_mac_out[8]_cal1_u149_mac ), .F2(dummy_abc_310_), .F3(dummy_abc_311_) );
      defparam ii1252.CONFIG_DATA = 16'h6666;
      defparam ii1252.PLACE_LOCATION = "NONE";
      defparam ii1252.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1253 ( .DX(nn1253), .F0(\a_mac_out[9]_cal1_u148_mac ), .F1(\a_mac_out[9]_cal1_u149_mac ), .F2(dummy_abc_312_), .F3(dummy_abc_313_) );
      defparam ii1253.CONFIG_DATA = 16'h6666;
      defparam ii1253.PLACE_LOCATION = "NONE";
      defparam ii1253.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1254 ( .DX(nn1254), .F0(\a_mac_out[10]_cal1_u148_mac ), .F1(\a_mac_out[10]_cal1_u149_mac ), .F2(dummy_abc_314_), .F3(dummy_abc_315_) );
      defparam ii1254.CONFIG_DATA = 16'h6666;
      defparam ii1254.PLACE_LOCATION = "NONE";
      defparam ii1254.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1255 ( .DX(nn1255), .F0(\a_mac_out[11]_cal1_u148_mac ), .F1(\a_mac_out[11]_cal1_u149_mac ), .F2(dummy_abc_316_), .F3(dummy_abc_317_) );
      defparam ii1255.CONFIG_DATA = 16'h6666;
      defparam ii1255.PLACE_LOCATION = "NONE";
      defparam ii1255.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1256 ( .DX(nn1256), .F0(\a_mac_out[12]_cal1_u148_mac ), .F1(\a_mac_out[12]_cal1_u149_mac ), .F2(dummy_abc_318_), .F3(dummy_abc_319_) );
      defparam ii1256.CONFIG_DATA = 16'h6666;
      defparam ii1256.PLACE_LOCATION = "NONE";
      defparam ii1256.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1257 ( .DX(nn1257), .F0(\a_mac_out[13]_cal1_u148_mac ), .F1(\a_mac_out[13]_cal1_u149_mac ), .F2(dummy_abc_320_), .F3(dummy_abc_321_) );
      defparam ii1257.CONFIG_DATA = 16'h6666;
      defparam ii1257.PLACE_LOCATION = "NONE";
      defparam ii1257.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1258 ( .DX(nn1258), .F0(dummy_abc_322_), .F1(dummy_abc_323_), .F2(dummy_abc_324_), .F3(dummy_abc_325_) );
      defparam ii1258.CONFIG_DATA = 16'h0000;
      defparam ii1258.PLACE_LOCATION = "NONE";
      defparam ii1258.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9_206_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u149_mac , 
              \a_mac_out[12]_cal1_u149_mac , \a_mac_out[11]_cal1_u149_mac , 
              \a_mac_out[10]_cal1_u149_mac , \a_mac_out[9]_cal1_u149_mac , \a_mac_out[8]_cal1_u149_mac , 
              \a_mac_out[7]_cal1_u149_mac , \a_mac_out[6]_cal1_u149_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_898_ ), 
        .DX( {nn1258, nn1257, nn1256, nn1255, nn1254, nn1253, nn1252, nn1251, 
              nn1250} ), 
        .SUM( {\cal1_u136_XORCI_SHIFT_0|SUM_net , 
              \cal1_u136_SUM_XORCI_0_151_|SUM_net , \cal1_u136_SUM_XORCI_0_148_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_145_|SUM_net , \cal1_u136_SUM_XORCI_0_142_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_139_|SUM_net , \cal1_u136_SUM_XORCI_0_136_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_133_|SUM_net , \cal1_u136_SUM_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1270 ( .DX(nn1270), .F0(\a_mac_out[6]_cal1_u146_mac ), .F1(\a_mac_out[6]_cal1_u147_mac ), .F2(nn1249), .F3(dummy_abc_326_) );
      defparam ii1270.CONFIG_DATA = 16'h9696;
      defparam ii1270.PLACE_LOCATION = "NONE";
      defparam ii1270.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1271 ( .DX(nn1271), .F0(\a_mac_out[6]_cal1_u146_mac ), .F1(\a_mac_out[6]_cal1_u147_mac ), .F2(dummy_abc_327_), .F3(dummy_abc_328_) );
      defparam ii1271.CONFIG_DATA = 16'h6666;
      defparam ii1271.PLACE_LOCATION = "NONE";
      defparam ii1271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1272 ( .DX(nn1272), .F0(\a_mac_out[7]_cal1_u146_mac ), .F1(\a_mac_out[7]_cal1_u147_mac ), .F2(dummy_abc_329_), .F3(dummy_abc_330_) );
      defparam ii1272.CONFIG_DATA = 16'h6666;
      defparam ii1272.PLACE_LOCATION = "NONE";
      defparam ii1272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1273 ( .DX(nn1273), .F0(\a_mac_out[8]_cal1_u146_mac ), .F1(\a_mac_out[8]_cal1_u147_mac ), .F2(dummy_abc_331_), .F3(dummy_abc_332_) );
      defparam ii1273.CONFIG_DATA = 16'h6666;
      defparam ii1273.PLACE_LOCATION = "NONE";
      defparam ii1273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1274 ( .DX(nn1274), .F0(\a_mac_out[9]_cal1_u146_mac ), .F1(\a_mac_out[9]_cal1_u147_mac ), .F2(dummy_abc_333_), .F3(dummy_abc_334_) );
      defparam ii1274.CONFIG_DATA = 16'h6666;
      defparam ii1274.PLACE_LOCATION = "NONE";
      defparam ii1274.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1275 ( .DX(nn1275), .F0(\a_mac_out[10]_cal1_u146_mac ), .F1(\a_mac_out[10]_cal1_u147_mac ), .F2(dummy_abc_335_), .F3(dummy_abc_336_) );
      defparam ii1275.CONFIG_DATA = 16'h6666;
      defparam ii1275.PLACE_LOCATION = "NONE";
      defparam ii1275.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1276 ( .DX(nn1276), .F0(\a_mac_out[11]_cal1_u146_mac ), .F1(\a_mac_out[11]_cal1_u147_mac ), .F2(dummy_abc_337_), .F3(dummy_abc_338_) );
      defparam ii1276.CONFIG_DATA = 16'h6666;
      defparam ii1276.PLACE_LOCATION = "NONE";
      defparam ii1276.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1277 ( .DX(nn1277), .F0(\a_mac_out[12]_cal1_u146_mac ), .F1(\a_mac_out[12]_cal1_u147_mac ), .F2(dummy_abc_339_), .F3(dummy_abc_340_) );
      defparam ii1277.CONFIG_DATA = 16'h6666;
      defparam ii1277.PLACE_LOCATION = "NONE";
      defparam ii1277.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1278 ( .DX(nn1278), .F0(\a_mac_out[13]_cal1_u146_mac ), .F1(\a_mac_out[13]_cal1_u147_mac ), .F2(dummy_abc_341_), .F3(dummy_abc_342_) );
      defparam ii1278.CONFIG_DATA = 16'h6666;
      defparam ii1278.PLACE_LOCATION = "NONE";
      defparam ii1278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1279 ( .DX(nn1279), .F0(dummy_abc_343_), .F1(dummy_abc_344_), .F2(dummy_abc_345_), .F3(dummy_abc_346_) );
      defparam ii1279.CONFIG_DATA = 16'h0000;
      defparam ii1279.PLACE_LOCATION = "NONE";
      defparam ii1279.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9_207_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u146_mac , 
              \a_mac_out[12]_cal1_u146_mac , \a_mac_out[11]_cal1_u146_mac , 
              \a_mac_out[10]_cal1_u146_mac , \a_mac_out[9]_cal1_u146_mac , \a_mac_out[8]_cal1_u146_mac , 
              \a_mac_out[7]_cal1_u146_mac , \a_mac_out[6]_cal1_u146_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_900_ ), 
        .DX( {nn1279, nn1278, nn1277, nn1276, nn1275, nn1274, nn1273, nn1272, 
              nn1271} ), 
        .SUM( {\cal1_u136_XORCI_SHIFT_1|SUM_net , 
              \cal1_u136_SUM_XORCI_1_172_|SUM_net , \cal1_u136_SUM_XORCI_1_169_|SUM_net , 
              \cal1_u136_SUM_XORCI_1_166_|SUM_net , \cal1_u136_SUM_XORCI_1_163_|SUM_net , 
              \cal1_u136_SUM_XORCI_1_160_|SUM_net , \cal1_u136_SUM_XORCI_1_157_|SUM_net , 
              \cal1_u136_SUM_XORCI_1_154_|SUM_net , \cal1_u136_SUM_XORCI_1|SUM_net } )
      );
    CS_LUT4_PRIM ii1291 ( .DX(nn1291), .F0(\cal1_u136_SUM_XORCI_0_133_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_154_|SUM_net ), .F2(dummy_abc_347_), .F3(dummy_abc_348_) );
      defparam ii1291.CONFIG_DATA = 16'h6666;
      defparam ii1291.PLACE_LOCATION = "NONE";
      defparam ii1291.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1292 ( .DX(nn1292), .F0(\cal1_u136_SUM_XORCI_0_136_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_157_|SUM_net ), .F2(dummy_abc_349_), .F3(dummy_abc_350_) );
      defparam ii1292.CONFIG_DATA = 16'h6666;
      defparam ii1292.PLACE_LOCATION = "NONE";
      defparam ii1292.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1293 ( .DX(nn1293), .F0(\cal1_u136_SUM_XORCI_0_139_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_160_|SUM_net ), .F2(dummy_abc_351_), .F3(dummy_abc_352_) );
      defparam ii1293.CONFIG_DATA = 16'h6666;
      defparam ii1293.PLACE_LOCATION = "NONE";
      defparam ii1293.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1294 ( .DX(nn1294), .F0(\cal1_u136_SUM_XORCI_0_142_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_163_|SUM_net ), .F2(dummy_abc_353_), .F3(dummy_abc_354_) );
      defparam ii1294.CONFIG_DATA = 16'h6666;
      defparam ii1294.PLACE_LOCATION = "NONE";
      defparam ii1294.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1295 ( .DX(nn1295), .F0(\cal1_u136_SUM_XORCI_0_145_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_166_|SUM_net ), .F2(dummy_abc_355_), .F3(dummy_abc_356_) );
      defparam ii1295.CONFIG_DATA = 16'h6666;
      defparam ii1295.PLACE_LOCATION = "NONE";
      defparam ii1295.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1296 ( .DX(nn1296), .F0(\cal1_u136_SUM_XORCI_0_148_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_169_|SUM_net ), .F2(dummy_abc_357_), .F3(dummy_abc_358_) );
      defparam ii1296.CONFIG_DATA = 16'h6666;
      defparam ii1296.PLACE_LOCATION = "NONE";
      defparam ii1296.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1297 ( .DX(nn1297), .F0(\cal1_u136_SUM_XORCI_0_151_|SUM_net ), .F1(\cal1_u136_SUM_XORCI_1_172_|SUM_net ), .F2(dummy_abc_359_), .F3(dummy_abc_360_) );
      defparam ii1297.CONFIG_DATA = 16'h6666;
      defparam ii1297.PLACE_LOCATION = "NONE";
      defparam ii1297.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1298 ( .DX(nn1298), .F0(dummy_abc_361_), .F1(dummy_abc_362_), .F2(dummy_abc_363_), .F3(dummy_abc_364_) );
      defparam ii1298.CONFIG_DATA = 16'h0000;
      defparam ii1298.PLACE_LOCATION = "NONE";
      defparam ii1298.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1299 ( .DX(nn1299), .F0(dummy_abc_365_), .F1(dummy_abc_366_), .F2(dummy_abc_367_), .F3(dummy_abc_368_) );
      defparam ii1299.CONFIG_DATA = 16'h0000;
      defparam ii1299.PLACE_LOCATION = "NONE";
      defparam ii1299.PCK_LOCATION = "NONE";
    scaler_ipc_adder_10 carry_10_208_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \cal1_u136_XORCI_SHIFT_0|SUM_net , 
              \cal1_u136_SUM_XORCI_0_151_|SUM_net , \cal1_u136_SUM_XORCI_0_148_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_145_|SUM_net , \cal1_u136_SUM_XORCI_0_142_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_139_|SUM_net , \cal1_u136_SUM_XORCI_0_136_|SUM_net , 
              \cal1_u136_SUM_XORCI_0_133_|SUM_net , nn1249} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_10_ ), 
        .DX( {nn1299, nn1298, nn1297, nn1296, nn1295, nn1294, nn1293, nn1292, 
              nn1291, nn1270} ), 
        .SUM( {dummy_11_, dummy_12_, dOut_7__net, dOut_6__net, dOut_5__net, 
              dOut_4__net, dOut_3__net, dOut_2__net, dOut_1__net, dOut_0__net} )
      );
    CS_LUT4_PRIM ii1312 ( .DX(nn1312), .F0(\a_mac_out[6]_cal1_u144_mac ), .F1(\a_mac_out[6]_cal1_u145_mac ), .F2(dummy_abc_369_), .F3(dummy_abc_370_) );
      defparam ii1312.CONFIG_DATA = 16'h6666;
      defparam ii1312.PLACE_LOCATION = "NONE";
      defparam ii1312.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1313 ( .DX(nn1313), .F0(\a_mac_out[6]_cal1_u144_mac ), .F1(\a_mac_out[6]_cal1_u145_mac ), .F2(dummy_abc_371_), .F3(dummy_abc_372_) );
      defparam ii1313.CONFIG_DATA = 16'h6666;
      defparam ii1313.PLACE_LOCATION = "NONE";
      defparam ii1313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1314 ( .DX(nn1314), .F0(\a_mac_out[7]_cal1_u144_mac ), .F1(\a_mac_out[7]_cal1_u145_mac ), .F2(dummy_abc_373_), .F3(dummy_abc_374_) );
      defparam ii1314.CONFIG_DATA = 16'h6666;
      defparam ii1314.PLACE_LOCATION = "NONE";
      defparam ii1314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1315 ( .DX(nn1315), .F0(\a_mac_out[8]_cal1_u144_mac ), .F1(\a_mac_out[8]_cal1_u145_mac ), .F2(dummy_abc_375_), .F3(dummy_abc_376_) );
      defparam ii1315.CONFIG_DATA = 16'h6666;
      defparam ii1315.PLACE_LOCATION = "NONE";
      defparam ii1315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1316 ( .DX(nn1316), .F0(\a_mac_out[9]_cal1_u144_mac ), .F1(\a_mac_out[9]_cal1_u145_mac ), .F2(dummy_abc_377_), .F3(dummy_abc_378_) );
      defparam ii1316.CONFIG_DATA = 16'h6666;
      defparam ii1316.PLACE_LOCATION = "NONE";
      defparam ii1316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1317 ( .DX(nn1317), .F0(\a_mac_out[10]_cal1_u144_mac ), .F1(\a_mac_out[10]_cal1_u145_mac ), .F2(dummy_abc_379_), .F3(dummy_abc_380_) );
      defparam ii1317.CONFIG_DATA = 16'h6666;
      defparam ii1317.PLACE_LOCATION = "NONE";
      defparam ii1317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1318 ( .DX(nn1318), .F0(\a_mac_out[11]_cal1_u144_mac ), .F1(\a_mac_out[11]_cal1_u145_mac ), .F2(dummy_abc_381_), .F3(dummy_abc_382_) );
      defparam ii1318.CONFIG_DATA = 16'h6666;
      defparam ii1318.PLACE_LOCATION = "NONE";
      defparam ii1318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1319 ( .DX(nn1319), .F0(\a_mac_out[12]_cal1_u144_mac ), .F1(\a_mac_out[12]_cal1_u145_mac ), .F2(dummy_abc_383_), .F3(dummy_abc_384_) );
      defparam ii1319.CONFIG_DATA = 16'h6666;
      defparam ii1319.PLACE_LOCATION = "NONE";
      defparam ii1319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1320 ( .DX(nn1320), .F0(\a_mac_out[13]_cal1_u144_mac ), .F1(\a_mac_out[13]_cal1_u145_mac ), .F2(dummy_abc_385_), .F3(dummy_abc_386_) );
      defparam ii1320.CONFIG_DATA = 16'h6666;
      defparam ii1320.PLACE_LOCATION = "NONE";
      defparam ii1320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1321 ( .DX(nn1321), .F0(dummy_abc_387_), .F1(dummy_abc_388_), .F2(dummy_abc_389_), .F3(dummy_abc_390_) );
      defparam ii1321.CONFIG_DATA = 16'h0000;
      defparam ii1321.PLACE_LOCATION = "NONE";
      defparam ii1321.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9_203_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u145_mac , 
              \a_mac_out[12]_cal1_u145_mac , \a_mac_out[11]_cal1_u145_mac , 
              \a_mac_out[10]_cal1_u145_mac , \a_mac_out[9]_cal1_u145_mac , \a_mac_out[8]_cal1_u145_mac , 
              \a_mac_out[7]_cal1_u145_mac , \a_mac_out[6]_cal1_u145_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_894_ ), 
        .DX( {nn1321, nn1320, nn1319, nn1318, nn1317, nn1316, nn1315, nn1314, 
              nn1313} ), 
        .SUM( {\cal1_u135_XORCI_SHIFT_0|SUM_net , 
              \cal1_u135_SUM_XORCI_0_85_|SUM_net , \cal1_u135_SUM_XORCI_0_82_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_79_|SUM_net , \cal1_u135_SUM_XORCI_0_76_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_73_|SUM_net , \cal1_u135_SUM_XORCI_0_70_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_67_|SUM_net , \cal1_u135_SUM_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1333 ( .DX(nn1333), .F0(\a_mac_out[6]_cal1_u142_mac ), .F1(\a_mac_out[6]_cal1_u143_mac ), .F2(nn1312), .F3(dummy_abc_391_) );
      defparam ii1333.CONFIG_DATA = 16'h9696;
      defparam ii1333.PLACE_LOCATION = "NONE";
      defparam ii1333.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1334 ( .DX(nn1334), .F0(\a_mac_out[6]_cal1_u142_mac ), .F1(\a_mac_out[6]_cal1_u143_mac ), .F2(dummy_abc_392_), .F3(dummy_abc_393_) );
      defparam ii1334.CONFIG_DATA = 16'h6666;
      defparam ii1334.PLACE_LOCATION = "NONE";
      defparam ii1334.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1335 ( .DX(nn1335), .F0(\a_mac_out[7]_cal1_u142_mac ), .F1(\a_mac_out[7]_cal1_u143_mac ), .F2(dummy_abc_394_), .F3(dummy_abc_395_) );
      defparam ii1335.CONFIG_DATA = 16'h6666;
      defparam ii1335.PLACE_LOCATION = "NONE";
      defparam ii1335.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1336 ( .DX(nn1336), .F0(\a_mac_out[8]_cal1_u142_mac ), .F1(\a_mac_out[8]_cal1_u143_mac ), .F2(dummy_abc_396_), .F3(dummy_abc_397_) );
      defparam ii1336.CONFIG_DATA = 16'h6666;
      defparam ii1336.PLACE_LOCATION = "NONE";
      defparam ii1336.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1337 ( .DX(nn1337), .F0(\a_mac_out[9]_cal1_u142_mac ), .F1(\a_mac_out[9]_cal1_u143_mac ), .F2(dummy_abc_398_), .F3(dummy_abc_399_) );
      defparam ii1337.CONFIG_DATA = 16'h6666;
      defparam ii1337.PLACE_LOCATION = "NONE";
      defparam ii1337.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1338 ( .DX(nn1338), .F0(\a_mac_out[10]_cal1_u142_mac ), .F1(\a_mac_out[10]_cal1_u143_mac ), .F2(dummy_abc_400_), .F3(dummy_abc_401_) );
      defparam ii1338.CONFIG_DATA = 16'h6666;
      defparam ii1338.PLACE_LOCATION = "NONE";
      defparam ii1338.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1339 ( .DX(nn1339), .F0(\a_mac_out[11]_cal1_u142_mac ), .F1(\a_mac_out[11]_cal1_u143_mac ), .F2(dummy_abc_402_), .F3(dummy_abc_403_) );
      defparam ii1339.CONFIG_DATA = 16'h6666;
      defparam ii1339.PLACE_LOCATION = "NONE";
      defparam ii1339.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1340 ( .DX(nn1340), .F0(\a_mac_out[12]_cal1_u142_mac ), .F1(\a_mac_out[12]_cal1_u143_mac ), .F2(dummy_abc_404_), .F3(dummy_abc_405_) );
      defparam ii1340.CONFIG_DATA = 16'h6666;
      defparam ii1340.PLACE_LOCATION = "NONE";
      defparam ii1340.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1341 ( .DX(nn1341), .F0(\a_mac_out[13]_cal1_u142_mac ), .F1(\a_mac_out[13]_cal1_u143_mac ), .F2(dummy_abc_406_), .F3(dummy_abc_407_) );
      defparam ii1341.CONFIG_DATA = 16'h6666;
      defparam ii1341.PLACE_LOCATION = "NONE";
      defparam ii1341.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1342 ( .DX(nn1342), .F0(dummy_abc_408_), .F1(dummy_abc_409_), .F2(dummy_abc_410_), .F3(dummy_abc_411_) );
      defparam ii1342.CONFIG_DATA = 16'h0000;
      defparam ii1342.PLACE_LOCATION = "NONE";
      defparam ii1342.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9_204_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u142_mac , 
              \a_mac_out[12]_cal1_u142_mac , \a_mac_out[11]_cal1_u142_mac , 
              \a_mac_out[10]_cal1_u142_mac , \a_mac_out[9]_cal1_u142_mac , \a_mac_out[8]_cal1_u142_mac , 
              \a_mac_out[7]_cal1_u142_mac , \a_mac_out[6]_cal1_u142_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_896_ ), 
        .DX( {nn1342, nn1341, nn1340, nn1339, nn1338, nn1337, nn1336, nn1335, 
              nn1334} ), 
        .SUM( {\cal1_u135_XORCI_SHIFT_1|SUM_net , 
              \cal1_u135_SUM_XORCI_1_106_|SUM_net , \cal1_u135_SUM_XORCI_1_103_|SUM_net , 
              \cal1_u135_SUM_XORCI_1_100_|SUM_net , \cal1_u135_SUM_XORCI_1_97_|SUM_net , 
              \cal1_u135_SUM_XORCI_1_94_|SUM_net , \cal1_u135_SUM_XORCI_1_91_|SUM_net , 
              \cal1_u135_SUM_XORCI_1_88_|SUM_net , \cal1_u135_SUM_XORCI_1|SUM_net } )
      );
    CS_LUT4_PRIM ii1354 ( .DX(nn1354), .F0(\cal1_u135_SUM_XORCI_0_67_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_88_|SUM_net ), .F2(dummy_abc_412_), .F3(dummy_abc_413_) );
      defparam ii1354.CONFIG_DATA = 16'h6666;
      defparam ii1354.PLACE_LOCATION = "NONE";
      defparam ii1354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1355 ( .DX(nn1355), .F0(\cal1_u135_SUM_XORCI_0_70_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_91_|SUM_net ), .F2(dummy_abc_414_), .F3(dummy_abc_415_) );
      defparam ii1355.CONFIG_DATA = 16'h6666;
      defparam ii1355.PLACE_LOCATION = "NONE";
      defparam ii1355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1356 ( .DX(nn1356), .F0(\cal1_u135_SUM_XORCI_0_73_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_94_|SUM_net ), .F2(dummy_abc_416_), .F3(dummy_abc_417_) );
      defparam ii1356.CONFIG_DATA = 16'h6666;
      defparam ii1356.PLACE_LOCATION = "NONE";
      defparam ii1356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1357 ( .DX(nn1357), .F0(\cal1_u135_SUM_XORCI_0_76_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_97_|SUM_net ), .F2(dummy_abc_418_), .F3(dummy_abc_419_) );
      defparam ii1357.CONFIG_DATA = 16'h6666;
      defparam ii1357.PLACE_LOCATION = "NONE";
      defparam ii1357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1358 ( .DX(nn1358), .F0(\cal1_u135_SUM_XORCI_0_79_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_100_|SUM_net ), .F2(dummy_abc_420_), .F3(dummy_abc_421_) );
      defparam ii1358.CONFIG_DATA = 16'h6666;
      defparam ii1358.PLACE_LOCATION = "NONE";
      defparam ii1358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1359 ( .DX(nn1359), .F0(\cal1_u135_SUM_XORCI_0_82_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_103_|SUM_net ), .F2(dummy_abc_422_), .F3(dummy_abc_423_) );
      defparam ii1359.CONFIG_DATA = 16'h6666;
      defparam ii1359.PLACE_LOCATION = "NONE";
      defparam ii1359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1360 ( .DX(nn1360), .F0(\cal1_u135_SUM_XORCI_0_85_|SUM_net ), .F1(\cal1_u135_SUM_XORCI_1_106_|SUM_net ), .F2(dummy_abc_424_), .F3(dummy_abc_425_) );
      defparam ii1360.CONFIG_DATA = 16'h6666;
      defparam ii1360.PLACE_LOCATION = "NONE";
      defparam ii1360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1361 ( .DX(nn1361), .F0(dummy_abc_426_), .F1(dummy_abc_427_), .F2(dummy_abc_428_), .F3(dummy_abc_429_) );
      defparam ii1361.CONFIG_DATA = 16'h0000;
      defparam ii1361.PLACE_LOCATION = "NONE";
      defparam ii1361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1362 ( .DX(nn1362), .F0(dummy_abc_430_), .F1(dummy_abc_431_), .F2(dummy_abc_432_), .F3(dummy_abc_433_) );
      defparam ii1362.CONFIG_DATA = 16'h0000;
      defparam ii1362.PLACE_LOCATION = "NONE";
      defparam ii1362.PCK_LOCATION = "NONE";
    scaler_ipc_adder_10 carry_10_205_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \cal1_u135_XORCI_SHIFT_0|SUM_net , 
              \cal1_u135_SUM_XORCI_0_85_|SUM_net , \cal1_u135_SUM_XORCI_0_82_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_79_|SUM_net , \cal1_u135_SUM_XORCI_0_76_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_73_|SUM_net , \cal1_u135_SUM_XORCI_0_70_|SUM_net , 
              \cal1_u135_SUM_XORCI_0_67_|SUM_net , nn1312} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_6_ ), 
        .DX( {nn1362, nn1361, nn1360, nn1359, nn1358, nn1357, nn1356, nn1355, 
              nn1354, nn1333} ), 
        .SUM( {dummy_7_, dummy_8_, dOut_15__net, dOut_14__net, dOut_13__net, 
              dOut_12__net, dOut_11__net, dOut_10__net, dOut_9__net, dOut_8__net} )
      );
    CS_LUT4_PRIM ii1375 ( .DX(nn1375), .F0(\a_mac_out[6]_cal1_u140_mac ), .F1(\a_mac_out[6]_cal1_u141_mac ), .F2(dummy_abc_434_), .F3(dummy_abc_435_) );
      defparam ii1375.CONFIG_DATA = 16'h6666;
      defparam ii1375.PLACE_LOCATION = "NONE";
      defparam ii1375.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1376 ( .DX(nn1376), .F0(\a_mac_out[6]_cal1_u140_mac ), .F1(\a_mac_out[6]_cal1_u141_mac ), .F2(dummy_abc_436_), .F3(dummy_abc_437_) );
      defparam ii1376.CONFIG_DATA = 16'h6666;
      defparam ii1376.PLACE_LOCATION = "NONE";
      defparam ii1376.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1377 ( .DX(nn1377), .F0(\a_mac_out[7]_cal1_u140_mac ), .F1(\a_mac_out[7]_cal1_u141_mac ), .F2(dummy_abc_438_), .F3(dummy_abc_439_) );
      defparam ii1377.CONFIG_DATA = 16'h6666;
      defparam ii1377.PLACE_LOCATION = "NONE";
      defparam ii1377.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1378 ( .DX(nn1378), .F0(\a_mac_out[8]_cal1_u140_mac ), .F1(\a_mac_out[8]_cal1_u141_mac ), .F2(dummy_abc_440_), .F3(dummy_abc_441_) );
      defparam ii1378.CONFIG_DATA = 16'h6666;
      defparam ii1378.PLACE_LOCATION = "NONE";
      defparam ii1378.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1379 ( .DX(nn1379), .F0(\a_mac_out[9]_cal1_u140_mac ), .F1(\a_mac_out[9]_cal1_u141_mac ), .F2(dummy_abc_442_), .F3(dummy_abc_443_) );
      defparam ii1379.CONFIG_DATA = 16'h6666;
      defparam ii1379.PLACE_LOCATION = "NONE";
      defparam ii1379.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1380 ( .DX(nn1380), .F0(\a_mac_out[10]_cal1_u140_mac ), .F1(\a_mac_out[10]_cal1_u141_mac ), .F2(dummy_abc_444_), .F3(dummy_abc_445_) );
      defparam ii1380.CONFIG_DATA = 16'h6666;
      defparam ii1380.PLACE_LOCATION = "NONE";
      defparam ii1380.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1381 ( .DX(nn1381), .F0(\a_mac_out[11]_cal1_u140_mac ), .F1(\a_mac_out[11]_cal1_u141_mac ), .F2(dummy_abc_446_), .F3(dummy_abc_447_) );
      defparam ii1381.CONFIG_DATA = 16'h6666;
      defparam ii1381.PLACE_LOCATION = "NONE";
      defparam ii1381.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1382 ( .DX(nn1382), .F0(\a_mac_out[12]_cal1_u140_mac ), .F1(\a_mac_out[12]_cal1_u141_mac ), .F2(dummy_abc_448_), .F3(dummy_abc_449_) );
      defparam ii1382.CONFIG_DATA = 16'h6666;
      defparam ii1382.PLACE_LOCATION = "NONE";
      defparam ii1382.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1383 ( .DX(nn1383), .F0(\a_mac_out[13]_cal1_u140_mac ), .F1(\a_mac_out[13]_cal1_u141_mac ), .F2(dummy_abc_450_), .F3(dummy_abc_451_) );
      defparam ii1383.CONFIG_DATA = 16'h6666;
      defparam ii1383.PLACE_LOCATION = "NONE";
      defparam ii1383.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1384 ( .DX(nn1384), .F0(dummy_abc_452_), .F1(dummy_abc_453_), .F2(dummy_abc_454_), .F3(dummy_abc_455_) );
      defparam ii1384.CONFIG_DATA = 16'h0000;
      defparam ii1384.PLACE_LOCATION = "NONE";
      defparam ii1384.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9 ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u141_mac , 
              \a_mac_out[12]_cal1_u141_mac , \a_mac_out[11]_cal1_u141_mac , 
              \a_mac_out[10]_cal1_u141_mac , \a_mac_out[9]_cal1_u141_mac , \a_mac_out[8]_cal1_u141_mac , 
              \a_mac_out[7]_cal1_u141_mac , \a_mac_out[6]_cal1_u141_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_890_ ), 
        .DX( {nn1384, nn1383, nn1382, nn1381, nn1380, nn1379, nn1378, nn1377, 
              nn1376} ), 
        .SUM( {\cal1_u134_XORCI_SHIFT_0|SUM_net , 
              \cal1_u134_SUM_XORCI_0_19_|SUM_net , \cal1_u134_SUM_XORCI_0_16_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_13_|SUM_net , \cal1_u134_SUM_XORCI_0_10_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_7_|SUM_net , \cal1_u134_SUM_XORCI_0_4_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_1_|SUM_net , \cal1_u134_SUM_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1396 ( .DX(nn1396), .F0(\a_mac_out[6]_cal1_u138_mac ), .F1(\a_mac_out[6]_cal1_u139_mac ), .F2(nn1375), .F3(dummy_abc_456_) );
      defparam ii1396.CONFIG_DATA = 16'h9696;
      defparam ii1396.PLACE_LOCATION = "NONE";
      defparam ii1396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1397 ( .DX(nn1397), .F0(\a_mac_out[6]_cal1_u138_mac ), .F1(\a_mac_out[6]_cal1_u139_mac ), .F2(dummy_abc_457_), .F3(dummy_abc_458_) );
      defparam ii1397.CONFIG_DATA = 16'h6666;
      defparam ii1397.PLACE_LOCATION = "NONE";
      defparam ii1397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1398 ( .DX(nn1398), .F0(\a_mac_out[7]_cal1_u138_mac ), .F1(\a_mac_out[7]_cal1_u139_mac ), .F2(dummy_abc_459_), .F3(dummy_abc_460_) );
      defparam ii1398.CONFIG_DATA = 16'h6666;
      defparam ii1398.PLACE_LOCATION = "NONE";
      defparam ii1398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1399 ( .DX(nn1399), .F0(\a_mac_out[8]_cal1_u138_mac ), .F1(\a_mac_out[8]_cal1_u139_mac ), .F2(dummy_abc_461_), .F3(dummy_abc_462_) );
      defparam ii1399.CONFIG_DATA = 16'h6666;
      defparam ii1399.PLACE_LOCATION = "NONE";
      defparam ii1399.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1400 ( .DX(nn1400), .F0(\a_mac_out[9]_cal1_u138_mac ), .F1(\a_mac_out[9]_cal1_u139_mac ), .F2(dummy_abc_463_), .F3(dummy_abc_464_) );
      defparam ii1400.CONFIG_DATA = 16'h6666;
      defparam ii1400.PLACE_LOCATION = "NONE";
      defparam ii1400.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1401 ( .DX(nn1401), .F0(\a_mac_out[10]_cal1_u138_mac ), .F1(\a_mac_out[10]_cal1_u139_mac ), .F2(dummy_abc_465_), .F3(dummy_abc_466_) );
      defparam ii1401.CONFIG_DATA = 16'h6666;
      defparam ii1401.PLACE_LOCATION = "NONE";
      defparam ii1401.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1402 ( .DX(nn1402), .F0(\a_mac_out[11]_cal1_u138_mac ), .F1(\a_mac_out[11]_cal1_u139_mac ), .F2(dummy_abc_467_), .F3(dummy_abc_468_) );
      defparam ii1402.CONFIG_DATA = 16'h6666;
      defparam ii1402.PLACE_LOCATION = "NONE";
      defparam ii1402.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1403 ( .DX(nn1403), .F0(\a_mac_out[12]_cal1_u138_mac ), .F1(\a_mac_out[12]_cal1_u139_mac ), .F2(dummy_abc_469_), .F3(dummy_abc_470_) );
      defparam ii1403.CONFIG_DATA = 16'h6666;
      defparam ii1403.PLACE_LOCATION = "NONE";
      defparam ii1403.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1404 ( .DX(nn1404), .F0(\a_mac_out[13]_cal1_u138_mac ), .F1(\a_mac_out[13]_cal1_u139_mac ), .F2(dummy_abc_471_), .F3(dummy_abc_472_) );
      defparam ii1404.CONFIG_DATA = 16'h6666;
      defparam ii1404.PLACE_LOCATION = "NONE";
      defparam ii1404.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1405 ( .DX(nn1405), .F0(dummy_abc_473_), .F1(dummy_abc_474_), .F2(dummy_abc_475_), .F3(dummy_abc_476_) );
      defparam ii1405.CONFIG_DATA = 16'h0000;
      defparam ii1405.PLACE_LOCATION = "NONE";
      defparam ii1405.PCK_LOCATION = "NONE";
    scaler_ipc_adder_9 carry_9_202_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[13]_cal1_u138_mac , 
              \a_mac_out[12]_cal1_u138_mac , \a_mac_out[11]_cal1_u138_mac , 
              \a_mac_out[10]_cal1_u138_mac , \a_mac_out[9]_cal1_u138_mac , \a_mac_out[8]_cal1_u138_mac , 
              \a_mac_out[7]_cal1_u138_mac , \a_mac_out[6]_cal1_u138_mac } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_892_ ), 
        .DX( {nn1405, nn1404, nn1403, nn1402, nn1401, nn1400, nn1399, nn1398, 
              nn1397} ), 
        .SUM( {\cal1_u134_XORCI_SHIFT_1|SUM_net , 
              \cal1_u134_SUM_XORCI_1_40_|SUM_net , \cal1_u134_SUM_XORCI_1_37_|SUM_net , 
              \cal1_u134_SUM_XORCI_1_34_|SUM_net , \cal1_u134_SUM_XORCI_1_31_|SUM_net , 
              \cal1_u134_SUM_XORCI_1_28_|SUM_net , \cal1_u134_SUM_XORCI_1_25_|SUM_net , 
              \cal1_u134_SUM_XORCI_1_22_|SUM_net , \cal1_u134_SUM_XORCI_1|SUM_net } )
      );
    CS_LUT4_PRIM ii1417 ( .DX(nn1417), .F0(\cal1_u134_SUM_XORCI_0_1_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_22_|SUM_net ), .F2(dummy_abc_477_), .F3(dummy_abc_478_) );
      defparam ii1417.CONFIG_DATA = 16'h6666;
      defparam ii1417.PLACE_LOCATION = "NONE";
      defparam ii1417.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1418 ( .DX(nn1418), .F0(\cal1_u134_SUM_XORCI_0_4_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_25_|SUM_net ), .F2(dummy_abc_479_), .F3(dummy_abc_480_) );
      defparam ii1418.CONFIG_DATA = 16'h6666;
      defparam ii1418.PLACE_LOCATION = "NONE";
      defparam ii1418.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1419 ( .DX(nn1419), .F0(\cal1_u134_SUM_XORCI_0_7_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_28_|SUM_net ), .F2(dummy_abc_481_), .F3(dummy_abc_482_) );
      defparam ii1419.CONFIG_DATA = 16'h6666;
      defparam ii1419.PLACE_LOCATION = "NONE";
      defparam ii1419.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1420 ( .DX(nn1420), .F0(\cal1_u134_SUM_XORCI_0_10_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_31_|SUM_net ), .F2(dummy_abc_483_), .F3(dummy_abc_484_) );
      defparam ii1420.CONFIG_DATA = 16'h6666;
      defparam ii1420.PLACE_LOCATION = "NONE";
      defparam ii1420.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1421 ( .DX(nn1421), .F0(\cal1_u134_SUM_XORCI_0_13_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_34_|SUM_net ), .F2(dummy_abc_485_), .F3(dummy_abc_486_) );
      defparam ii1421.CONFIG_DATA = 16'h6666;
      defparam ii1421.PLACE_LOCATION = "NONE";
      defparam ii1421.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1422 ( .DX(nn1422), .F0(\cal1_u134_SUM_XORCI_0_16_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_37_|SUM_net ), .F2(dummy_abc_487_), .F3(dummy_abc_488_) );
      defparam ii1422.CONFIG_DATA = 16'h6666;
      defparam ii1422.PLACE_LOCATION = "NONE";
      defparam ii1422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1423 ( .DX(nn1423), .F0(\cal1_u134_SUM_XORCI_0_19_|SUM_net ), .F1(\cal1_u134_SUM_XORCI_1_40_|SUM_net ), .F2(dummy_abc_489_), .F3(dummy_abc_490_) );
      defparam ii1423.CONFIG_DATA = 16'h6666;
      defparam ii1423.PLACE_LOCATION = "NONE";
      defparam ii1423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1424 ( .DX(nn1424), .F0(dummy_abc_491_), .F1(dummy_abc_492_), .F2(dummy_abc_493_), .F3(dummy_abc_494_) );
      defparam ii1424.CONFIG_DATA = 16'h0000;
      defparam ii1424.PLACE_LOCATION = "NONE";
      defparam ii1424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1425 ( .DX(nn1425), .F0(dummy_abc_495_), .F1(dummy_abc_496_), .F2(dummy_abc_497_), .F3(dummy_abc_498_) );
      defparam ii1425.CONFIG_DATA = 16'h0000;
      defparam ii1425.PLACE_LOCATION = "NONE";
      defparam ii1425.PCK_LOCATION = "NONE";
    scaler_ipc_adder_10 carry_10 ( 
        .CA( {a_acc_en_cal1_u137_mac, \cal1_u134_XORCI_SHIFT_0|SUM_net , 
              \cal1_u134_SUM_XORCI_0_19_|SUM_net , \cal1_u134_SUM_XORCI_0_16_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_13_|SUM_net , \cal1_u134_SUM_XORCI_0_10_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_7_|SUM_net , \cal1_u134_SUM_XORCI_0_4_|SUM_net , 
              \cal1_u134_SUM_XORCI_0_1_|SUM_net , nn1375} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_2_ ), 
        .DX( {nn1425, nn1424, nn1423, nn1422, nn1421, nn1420, nn1419, nn1418, 
              nn1417, nn1396} ), 
        .SUM( {dummy_3_, dummy_4_, dOut_23__net, dOut_22__net, dOut_21__net, 
              dOut_20__net, dOut_19__net, dOut_18__net, dOut_17__net, dOut_16__net} )
      );
    CS_LUT4_PRIM ii1438 ( .DX(nn1438), .F0(outYRes[0]), .F1(\cal1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_499_), .F3(dummy_abc_500_) );
      defparam ii1438.CONFIG_DATA = 16'h9999;
      defparam ii1438.PLACE_LOCATION = "NONE";
      defparam ii1438.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1439 ( .DX(nn1439), .F0(outYRes[1]), .F1(\cal1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_501_), .F3(dummy_abc_502_) );
      defparam ii1439.CONFIG_DATA = 16'h9999;
      defparam ii1439.PLACE_LOCATION = "NONE";
      defparam ii1439.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1440 ( .DX(nn1440), .F0(outYRes[2]), .F1(\cal1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_503_), .F3(dummy_abc_504_) );
      defparam ii1440.CONFIG_DATA = 16'h9999;
      defparam ii1440.PLACE_LOCATION = "NONE";
      defparam ii1440.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1441 ( .DX(nn1441), .F0(outYRes[3]), .F1(\cal1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_505_), .F3(dummy_abc_506_) );
      defparam ii1441.CONFIG_DATA = 16'h9999;
      defparam ii1441.PLACE_LOCATION = "NONE";
      defparam ii1441.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1442 ( .DX(nn1442), .F0(outYRes[4]), .F1(\cal1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_507_), .F3(dummy_abc_508_) );
      defparam ii1442.CONFIG_DATA = 16'h9999;
      defparam ii1442.PLACE_LOCATION = "NONE";
      defparam ii1442.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1443 ( .DX(nn1443), .F0(outYRes[5]), .F1(\cal1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_509_), .F3(dummy_abc_510_) );
      defparam ii1443.CONFIG_DATA = 16'h9999;
      defparam ii1443.PLACE_LOCATION = "NONE";
      defparam ii1443.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1444 ( .DX(nn1444), .F0(outYRes[6]), .F1(\cal1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_511_), .F3(dummy_abc_512_) );
      defparam ii1444.CONFIG_DATA = 16'h9999;
      defparam ii1444.PLACE_LOCATION = "NONE";
      defparam ii1444.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1445 ( .DX(nn1445), .F0(outYRes[7]), .F1(\cal1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_513_), .F3(dummy_abc_514_) );
      defparam ii1445.CONFIG_DATA = 16'h9999;
      defparam ii1445.PLACE_LOCATION = "NONE";
      defparam ii1445.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1446 ( .DX(nn1446), .F0(outYRes[8]), .F1(\cal1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_515_), .F3(dummy_abc_516_) );
      defparam ii1446.CONFIG_DATA = 16'h9999;
      defparam ii1446.PLACE_LOCATION = "NONE";
      defparam ii1446.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1447 ( .DX(nn1447), .F0(outYRes[9]), .F1(\cal1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_517_), .F3(dummy_abc_518_) );
      defparam ii1447.CONFIG_DATA = 16'h9999;
      defparam ii1447.PLACE_LOCATION = "NONE";
      defparam ii1447.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1448 ( .DX(nn1448), .F0(outYRes[10]), .F1(\cal1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_519_), .F3(dummy_abc_520_) );
      defparam ii1448.CONFIG_DATA = 16'h9999;
      defparam ii1448.PLACE_LOCATION = "NONE";
      defparam ii1448.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1449 ( .DX(nn1449), .F0(dummy_abc_521_), .F1(dummy_abc_522_), .F2(dummy_abc_523_), .F3(dummy_abc_524_) );
      defparam ii1449.CONFIG_DATA = 16'hFFFF;
      defparam ii1449.PLACE_LOCATION = "NONE";
      defparam ii1449.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_211_ ( 
        .CA( {a_acc_en_cal1_u137_mac, outYRes[10], outYRes[9], outYRes[8], 
              outYRes[7], outYRes[6], outYRes[5], outYRes[4], outYRes[3], outYRes[2], 
              outYRes[1], outYRes[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_36_ ), 
        .DX( {nn1449, nn1448, nn1447, nn1446, nn1445, nn1444, nn1443, nn1442, 
              nn1441, nn1440, nn1439, nn1438} ), 
        .SUM( {\cal1_u59_XORCI_11|SUM_net , dummy_37_, dummy_38_, dummy_39_, 
              dummy_40_, dummy_41_, dummy_42_, dummy_43_, dummy_44_, dummy_45_, 
              dummy_46_, dummy_47_} )
      );
    CS_LUT4_PRIM ii1464 ( .DX(nn1464), .F0(outXRes[0]), .F1(\cal1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_525_), .F3(dummy_abc_526_) );
      defparam ii1464.CONFIG_DATA = 16'h9999;
      defparam ii1464.PLACE_LOCATION = "NONE";
      defparam ii1464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1465 ( .DX(nn1465), .F0(outXRes[1]), .F1(\cal1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_527_), .F3(dummy_abc_528_) );
      defparam ii1465.CONFIG_DATA = 16'h9999;
      defparam ii1465.PLACE_LOCATION = "NONE";
      defparam ii1465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1466 ( .DX(nn1466), .F0(outXRes[2]), .F1(\cal1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_529_), .F3(dummy_abc_530_) );
      defparam ii1466.CONFIG_DATA = 16'h9999;
      defparam ii1466.PLACE_LOCATION = "NONE";
      defparam ii1466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1467 ( .DX(nn1467), .F0(outXRes[3]), .F1(\cal1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_531_), .F3(dummy_abc_532_) );
      defparam ii1467.CONFIG_DATA = 16'h9999;
      defparam ii1467.PLACE_LOCATION = "NONE";
      defparam ii1467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1468 ( .DX(nn1468), .F0(outXRes[4]), .F1(\cal1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_533_), .F3(dummy_abc_534_) );
      defparam ii1468.CONFIG_DATA = 16'h9999;
      defparam ii1468.PLACE_LOCATION = "NONE";
      defparam ii1468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1469 ( .DX(nn1469), .F0(outXRes[5]), .F1(\cal1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_535_), .F3(dummy_abc_536_) );
      defparam ii1469.CONFIG_DATA = 16'h9999;
      defparam ii1469.PLACE_LOCATION = "NONE";
      defparam ii1469.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1470 ( .DX(nn1470), .F0(outXRes[6]), .F1(\cal1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_537_), .F3(dummy_abc_538_) );
      defparam ii1470.CONFIG_DATA = 16'h9999;
      defparam ii1470.PLACE_LOCATION = "NONE";
      defparam ii1470.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1471 ( .DX(nn1471), .F0(outXRes[7]), .F1(\cal1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_539_), .F3(dummy_abc_540_) );
      defparam ii1471.CONFIG_DATA = 16'h9999;
      defparam ii1471.PLACE_LOCATION = "NONE";
      defparam ii1471.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1472 ( .DX(nn1472), .F0(outXRes[8]), .F1(\cal1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_541_), .F3(dummy_abc_542_) );
      defparam ii1472.CONFIG_DATA = 16'h9999;
      defparam ii1472.PLACE_LOCATION = "NONE";
      defparam ii1472.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1473 ( .DX(nn1473), .F0(outXRes[9]), .F1(\cal1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_543_), .F3(dummy_abc_544_) );
      defparam ii1473.CONFIG_DATA = 16'h9999;
      defparam ii1473.PLACE_LOCATION = "NONE";
      defparam ii1473.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1474 ( .DX(nn1474), .F0(outXRes[10]), .F1(\cal1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_545_), .F3(dummy_abc_546_) );
      defparam ii1474.CONFIG_DATA = 16'h9999;
      defparam ii1474.PLACE_LOCATION = "NONE";
      defparam ii1474.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1475 ( .DX(nn1475), .F0(dummy_abc_547_), .F1(dummy_abc_548_), .F2(dummy_abc_549_), .F3(dummy_abc_550_) );
      defparam ii1475.CONFIG_DATA = 16'hFFFF;
      defparam ii1475.PLACE_LOCATION = "NONE";
      defparam ii1475.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12 ( 
        .CA( {a_acc_en_cal1_u137_mac, outXRes[10], outXRes[9], outXRes[8], 
              outXRes[7], outXRes[6], outXRes[5], outXRes[4], outXRes[3], outXRes[2], 
              outXRes[1], outXRes[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_23_ ), 
        .DX( {nn1475, nn1474, nn1473, nn1472, nn1471, nn1470, nn1469, nn1468, 
              nn1467, nn1466, nn1465, nn1464} ), 
        .SUM( {\cal1_u57_XORCI_11|SUM_net , dummy_24_, dummy_25_, dummy_26_, 
              dummy_27_, dummy_28_, dummy_29_, dummy_30_, dummy_31_, dummy_32_, 
              dummy_33_, dummy_34_} )
      );
    CS_LUT4_PRIM ii1490 ( .DX(nn1490), .F0(\cal1_enforceJmp__reg|Q_net ), .F1(\cal1_jmp1Normal__reg|Q_net ), .F2(dummy_abc_551_), .F3(dummy_abc_552_) );
      defparam ii1490.CONFIG_DATA = 16'h1111;
      defparam ii1490.PLACE_LOCATION = "NONE";
      defparam ii1490.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1491 ( .DX(u8218_Y), .F0(rst), .F1(u8245_IN), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(nn1490) );
      defparam ii1491.CONFIG_DATA = 16'h1441;
      defparam ii1491.PLACE_LOCATION = "NONE";
      defparam ii1491.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1492 ( .DX(nn1492), .F0(u8245_D0), .F1(u8245_I0_3_), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(u8218_Y) );
      defparam ii1492.CONFIG_DATA = 16'h3ACA;
      defparam ii1492.PLACE_LOCATION = "NONE";
      defparam ii1492.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1493 ( .DX(nn1493), .F0(u8245_I0), .F1(u8245_I0_0_), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(u8218_Y) );
      defparam ii1493.CONFIG_DATA = 16'h5553;
      defparam ii1493.PLACE_LOCATION = "NONE";
      defparam ii1493.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1494 ( .DX(nn1494), .F0(\cal1_jmp2Normal__reg|Q_net ), .F1(nn1490), .F2(nn1492), .F3(nn1493) );
      defparam ii1494.CONFIG_DATA = 16'h8CBF;
      defparam ii1494.PLACE_LOCATION = "NONE";
      defparam ii1494.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1495 ( .DX(nn1495), .F0(rst), .F1(u8245_I0_0_), .F2(nn1490), .F3(dummy_abc_553_) );
      defparam ii1495.CONFIG_DATA = 16'h1010;
      defparam ii1495.PLACE_LOCATION = "NONE";
      defparam ii1495.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1496 ( .DX(nn1496), .F0(u8245_I0), .F1(\inputctrl1_jmp__reg|Q_net ), .F2(u8218_Y), .F3(nn1495) );
      defparam ii1496.CONFIG_DATA = 16'h7F40;
      defparam ii1496.PLACE_LOCATION = "NONE";
      defparam ii1496.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1497 ( .DX(u5018_OUT), .F0(rst), .F1(\cal1_jmp2Normal__reg|Q_net ), .F2(nn1494), .F3(nn1496) );
      defparam ii1497.CONFIG_DATA = 16'h32FA;
      defparam ii1497.PLACE_LOCATION = "NONE";
      defparam ii1497.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1498 ( .DX(nn1498), .F0(HS_2079_net), .F1(\cal1_VSNormal__reg|Q_net ), .F2(\cal1_enforceJmp__reg|Q_net ), .F3(dummy_abc_554_) );
      defparam ii1498.CONFIG_DATA = 16'h0101;
      defparam ii1498.PLACE_LOCATION = "NONE";
      defparam ii1498.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1499 ( .DX(nn1499), .F0(u8245_IN), .F1(dummy_62_), .F2(u5018_OUT), .F3(nn1498) );
      defparam ii1499.CONFIG_DATA = 16'h8F00;
      defparam ii1499.PLACE_LOCATION = "NONE";
      defparam ii1499.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1500 ( .DX(nn1500), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(\cal1_xAddress__reg[3]|Q_net ), .F2(\cal1_xAddress__reg[4]|Q_net ), .F3(\cal1_xAddress__reg[5]|Q_net ) );
      defparam ii1500.CONFIG_DATA = 16'h0001;
      defparam ii1500.PLACE_LOCATION = "NONE";
      defparam ii1500.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1501 ( .DX(nn1501), .F0(\cal1_xAddress__reg[10]|Q_net ), .F1(\cal1_xAddress__reg[1]|Q_net ), .F2(\cal1_xAddress__reg[6]|Q_net ), .F3(nn1500) );
      defparam ii1501.CONFIG_DATA = 16'h0100;
      defparam ii1501.PLACE_LOCATION = "NONE";
      defparam ii1501.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1502 ( .DX(nn1502), .F0(\cal1_xAddress__reg[7]|Q_net ), .F1(\cal1_xAddress__reg[8]|Q_net ), .F2(\cal1_xAddress__reg[9]|Q_net ), .F3(nn1501) );
      defparam ii1502.CONFIG_DATA = 16'h0100;
      defparam ii1502.PLACE_LOCATION = "NONE";
      defparam ii1502.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1503 ( .DX(nn1503), .F0(\cal1_yAddress__reg[3]|Q_net ), .F1(\cal1_yAddress__reg[4]|Q_net ), .F2(\cal1_yAddress__reg[5]|Q_net ), .F3(\cal1_yAddress__reg[6]|Q_net ) );
      defparam ii1503.CONFIG_DATA = 16'h0001;
      defparam ii1503.PLACE_LOCATION = "NONE";
      defparam ii1503.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1504 ( .DX(nn1504), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(\cal1_yAddress__reg[10]|Q_net ), .F2(\cal1_yAddress__reg[1]|Q_net ), .F3(nn1503) );
      defparam ii1504.CONFIG_DATA = 16'h0100;
      defparam ii1504.PLACE_LOCATION = "NONE";
      defparam ii1504.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1505 ( .DX(nn1505), .F0(\cal1_yAddress__reg[7]|Q_net ), .F1(\cal1_yAddress__reg[8]|Q_net ), .F2(\cal1_yAddress__reg[9]|Q_net ), .F3(nn1504) );
      defparam ii1505.CONFIG_DATA = 16'h0100;
      defparam ii1505.PLACE_LOCATION = "NONE";
      defparam ii1505.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1506 ( .DX(nn1506), .F0(\cal1_xAddress__reg[2]|Q_net ), .F1(\cal1_yAddress__reg[2]|Q_net ), .F2(nn1502), .F3(nn1505) );
      defparam ii1506.CONFIG_DATA = 16'h8CAF;
      defparam ii1506.PLACE_LOCATION = "NONE";
      defparam ii1506.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1507 ( .DX(dOutEn), .F0(dummy_36_), .F1(dummy_23_), .F2(nn1499), .F3(nn1506) );
      defparam ii1507.CONFIG_DATA = 16'h8000;
      defparam ii1507.PLACE_LOCATION = "NONE";
      defparam ii1507.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1508 ( .DX(\haa[0]_fifo1_ram_inst_0A_u_emb18k_0 ), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F2(u8231_O), .F3(dummy_abc_555_) );
      defparam ii1508.CONFIG_DATA = 16'hCACA;
      defparam ii1508.PLACE_LOCATION = "NONE";
      defparam ii1508.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1509 ( .DX(\haa[0]_fifo1_ram_inst_1A_u_emb18k_0 ), .F0(rst), .F1(\cal1_ramRdAddr__reg[10]|Q_net ), .F2(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F3(u8231_O) );
      defparam ii1509.CONFIG_DATA = 16'hD8CC;
      defparam ii1509.PLACE_LOCATION = "NONE";
      defparam ii1509.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1510 ( .DX(u8205_O), .F0(u5018_OUT), .F1(dummy_abc_556_), .F2(dummy_abc_557_), .F3(dummy_abc_558_) );
      defparam ii1510.CONFIG_DATA = 16'h5555;
      defparam ii1510.PLACE_LOCATION = "NONE";
      defparam ii1510.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1511 ( .DX(nn1511), .F0(\cal1_jmp2Normal__reg|Q_net ), .F1(nn1490), .F2(dummy_abc_559_), .F3(dummy_abc_560_) );
      defparam ii1511.CONFIG_DATA = 16'h8888;
      defparam ii1511.PLACE_LOCATION = "NONE";
      defparam ii1511.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1512 ( .DX(nn1512), .F0(u5502_I1_5_), .F1(nn1490), .F2(dummy_abc_561_), .F3(dummy_abc_562_) );
      defparam ii1512.CONFIG_DATA = 16'h2222;
      defparam ii1512.PLACE_LOCATION = "NONE";
      defparam ii1512.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1513 ( .DX(u8224_O), .F0(rst), .F1(u5502_I1), .F2(nn1511), .F3(nn1512) );
      defparam ii1513.CONFIG_DATA = 16'hFFEA;
      defparam ii1513.PLACE_LOCATION = "NONE";
      defparam ii1513.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1514 ( .DX(u8230_O), .F0(rst), .F1(u5502_IN), .F2(nn1511), .F3(nn1512) );
      defparam ii1514.CONFIG_DATA = 16'h5540;
      defparam ii1514.PLACE_LOCATION = "NONE";
      defparam ii1514.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1515 ( .DX(wea_fifo1_ram_inst_0A_u_emb18k_0), .F0(rst), .F1(u5859_I1), .F2(\inputctrl1_jmp__reg|Q_net ), .F3(\inputctrl1_ramWrtEn__reg|Q_net ) );
      defparam ii1515.CONFIG_DATA = 16'hEA00;
      defparam ii1515.PLACE_LOCATION = "NONE";
      defparam ii1515.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1516 ( .DX(wea_fifo1_ram_inst_1A_u_emb18k_0), .F0(rst), .F1(\inputctrl1_ramWrtEn__reg|Q_net ), .F2(u8231_O), .F3(dummy_abc_563_) );
      defparam ii1516.CONFIG_DATA = 16'h4040;
      defparam ii1516.PLACE_LOCATION = "NONE";
      defparam ii1516.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1517 ( .DX(nn1517), .F0(dummy_36_), .F1(dummy_23_), .F2(dummy_abc_564_), .F3(dummy_abc_565_) );
      defparam ii1517.CONFIG_DATA = 16'h2222;
      defparam ii1517.PLACE_LOCATION = "NONE";
      defparam ii1517.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1518 ( .DX(nn1518), .F0(dummy_36_), .F1(dummy_23_), .F2(dummy_abc_566_), .F3(dummy_abc_567_) );
      defparam ii1518.CONFIG_DATA = 16'h7777;
      defparam ii1518.PLACE_LOCATION = "NONE";
      defparam ii1518.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1519 ( .DX(nn1519), .F0(\cal1_VSNormal__reg|Q_net ), .F1(dummy_36_), .F2(nn1518), .F3(dummy_abc_568_) );
      defparam ii1519.CONFIG_DATA = 16'hB0B0;
      defparam ii1519.PLACE_LOCATION = "NONE";
      defparam ii1519.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1520 ( .DX(nn1520), .F0(\cal1_jmp1Normal__reg|Q_net ), .F1(dummy_62_), .F2(dummy_abc_569_), .F3(dummy_abc_570_) );
      defparam ii1520.CONFIG_DATA = 16'h1111;
      defparam ii1520.PLACE_LOCATION = "NONE";
      defparam ii1520.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1521 ( .DX(nn1521), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_571_), .F3(dummy_abc_572_) );
      defparam ii1521.CONFIG_DATA = 16'h9999;
      defparam ii1521.PLACE_LOCATION = "NONE";
      defparam ii1521.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1522 ( .DX(nn1522), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_573_), .F3(dummy_abc_574_) );
      defparam ii1522.CONFIG_DATA = 16'h9999;
      defparam ii1522.PLACE_LOCATION = "NONE";
      defparam ii1522.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1523 ( .DX(nn1523), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_abc_575_), .F3(dummy_abc_576_) );
      defparam ii1523.CONFIG_DATA = 16'h9999;
      defparam ii1523.PLACE_LOCATION = "NONE";
      defparam ii1523.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1524 ( .DX(nn1524), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[3]|Q_net ), .F2(dummy_abc_577_), .F3(dummy_abc_578_) );
      defparam ii1524.CONFIG_DATA = 16'h9999;
      defparam ii1524.PLACE_LOCATION = "NONE";
      defparam ii1524.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1525 ( .DX(nn1525), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[4]|Q_net ), .F2(dummy_abc_579_), .F3(dummy_abc_580_) );
      defparam ii1525.CONFIG_DATA = 16'h9999;
      defparam ii1525.PLACE_LOCATION = "NONE";
      defparam ii1525.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1526 ( .DX(nn1526), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[5]|Q_net ), .F2(dummy_abc_581_), .F3(dummy_abc_582_) );
      defparam ii1526.CONFIG_DATA = 16'h9999;
      defparam ii1526.PLACE_LOCATION = "NONE";
      defparam ii1526.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1527 ( .DX(nn1527), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[6]|Q_net ), .F2(dummy_abc_583_), .F3(dummy_abc_584_) );
      defparam ii1527.CONFIG_DATA = 16'h9999;
      defparam ii1527.PLACE_LOCATION = "NONE";
      defparam ii1527.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1528 ( .DX(nn1528), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[7]|Q_net ), .F2(dummy_abc_585_), .F3(dummy_abc_586_) );
      defparam ii1528.CONFIG_DATA = 16'h9999;
      defparam ii1528.PLACE_LOCATION = "NONE";
      defparam ii1528.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1529 ( .DX(nn1529), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[8]|Q_net ), .F2(dummy_abc_587_), .F3(dummy_abc_588_) );
      defparam ii1529.CONFIG_DATA = 16'h9999;
      defparam ii1529.PLACE_LOCATION = "NONE";
      defparam ii1529.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1530 ( .DX(nn1530), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[9]|Q_net ), .F2(dummy_abc_589_), .F3(dummy_abc_590_) );
      defparam ii1530.CONFIG_DATA = 16'h9999;
      defparam ii1530.PLACE_LOCATION = "NONE";
      defparam ii1530.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1531 ( .DX(nn1531), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[10]|Q_net ), .F2(dummy_abc_591_), .F3(dummy_abc_592_) );
      defparam ii1531.CONFIG_DATA = 16'h9999;
      defparam ii1531.PLACE_LOCATION = "NONE";
      defparam ii1531.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1532 ( .DX(nn1532), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[11]|Q_net ), .F2(dummy_abc_593_), .F3(dummy_abc_594_) );
      defparam ii1532.CONFIG_DATA = 16'h9999;
      defparam ii1532.PLACE_LOCATION = "NONE";
      defparam ii1532.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1533 ( .DX(nn1533), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[12]|Q_net ), .F2(dummy_abc_595_), .F3(dummy_abc_596_) );
      defparam ii1533.CONFIG_DATA = 16'h9999;
      defparam ii1533.PLACE_LOCATION = "NONE";
      defparam ii1533.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1534 ( .DX(nn1534), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[13]|Q_net ), .F2(dummy_abc_597_), .F3(dummy_abc_598_) );
      defparam ii1534.CONFIG_DATA = 16'h9999;
      defparam ii1534.PLACE_LOCATION = "NONE";
      defparam ii1534.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1535 ( .DX(nn1535), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[14]|Q_net ), .F2(dummy_abc_599_), .F3(dummy_abc_600_) );
      defparam ii1535.CONFIG_DATA = 16'h9999;
      defparam ii1535.PLACE_LOCATION = "NONE";
      defparam ii1535.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1536 ( .DX(nn1536), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[15]|Q_net ), .F2(dummy_abc_601_), .F3(dummy_abc_602_) );
      defparam ii1536.CONFIG_DATA = 16'h9999;
      defparam ii1536.PLACE_LOCATION = "NONE";
      defparam ii1536.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1537 ( .DX(nn1537), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_603_), .F3(dummy_abc_604_) );
      defparam ii1537.CONFIG_DATA = 16'h9999;
      defparam ii1537.PLACE_LOCATION = "NONE";
      defparam ii1537.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1538 ( .DX(nn1538), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_605_), .F3(dummy_abc_606_) );
      defparam ii1538.CONFIG_DATA = 16'h9999;
      defparam ii1538.PLACE_LOCATION = "NONE";
      defparam ii1538.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1539 ( .DX(nn1539), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_abc_607_), .F2(dummy_abc_608_), .F3(dummy_abc_609_) );
      defparam ii1539.CONFIG_DATA = 16'h5555;
      defparam ii1539.PLACE_LOCATION = "NONE";
      defparam ii1539.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1540 ( .DX(nn1540), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_610_), .F2(dummy_abc_611_), .F3(dummy_abc_612_) );
      defparam ii1540.CONFIG_DATA = 16'h5555;
      defparam ii1540.PLACE_LOCATION = "NONE";
      defparam ii1540.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1541 ( .DX(nn1541), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_613_), .F2(dummy_abc_614_), .F3(dummy_abc_615_) );
      defparam ii1541.CONFIG_DATA = 16'h5555;
      defparam ii1541.PLACE_LOCATION = "NONE";
      defparam ii1541.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1542 ( .DX(nn1542), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_616_), .F2(dummy_abc_617_), .F3(dummy_abc_618_) );
      defparam ii1542.CONFIG_DATA = 16'h5555;
      defparam ii1542.PLACE_LOCATION = "NONE";
      defparam ii1542.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1543 ( .DX(nn1543), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_619_), .F2(dummy_abc_620_), .F3(dummy_abc_621_) );
      defparam ii1543.CONFIG_DATA = 16'h5555;
      defparam ii1543.PLACE_LOCATION = "NONE";
      defparam ii1543.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1544 ( .DX(nn1544), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_622_), .F2(dummy_abc_623_), .F3(dummy_abc_624_) );
      defparam ii1544.CONFIG_DATA = 16'h5555;
      defparam ii1544.PLACE_LOCATION = "NONE";
      defparam ii1544.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1545 ( .DX(nn1545), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_625_), .F2(dummy_abc_626_), .F3(dummy_abc_627_) );
      defparam ii1545.CONFIG_DATA = 16'h5555;
      defparam ii1545.PLACE_LOCATION = "NONE";
      defparam ii1545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1546 ( .DX(nn1546), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_628_), .F2(dummy_abc_629_), .F3(dummy_abc_630_) );
      defparam ii1546.CONFIG_DATA = 16'h5555;
      defparam ii1546.PLACE_LOCATION = "NONE";
      defparam ii1546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1547 ( .DX(nn1547), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_631_), .F2(dummy_abc_632_), .F3(dummy_abc_633_) );
      defparam ii1547.CONFIG_DATA = 16'h5555;
      defparam ii1547.PLACE_LOCATION = "NONE";
      defparam ii1547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1548 ( .DX(nn1548), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_634_), .F2(dummy_abc_635_), .F3(dummy_abc_636_) );
      defparam ii1548.CONFIG_DATA = 16'h5555;
      defparam ii1548.PLACE_LOCATION = "NONE";
      defparam ii1548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1549 ( .DX(nn1549), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_637_), .F2(dummy_abc_638_), .F3(dummy_abc_639_) );
      defparam ii1549.CONFIG_DATA = 16'h5555;
      defparam ii1549.PLACE_LOCATION = "NONE";
      defparam ii1549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1550 ( .DX(nn1550), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_640_), .F2(dummy_abc_641_), .F3(dummy_abc_642_) );
      defparam ii1550.CONFIG_DATA = 16'h5555;
      defparam ii1550.PLACE_LOCATION = "NONE";
      defparam ii1550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1551 ( .DX(nn1551), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_643_), .F2(dummy_abc_644_), .F3(dummy_abc_645_) );
      defparam ii1551.CONFIG_DATA = 16'h5555;
      defparam ii1551.PLACE_LOCATION = "NONE";
      defparam ii1551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1552 ( .DX(nn1552), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_646_), .F2(dummy_abc_647_), .F3(dummy_abc_648_) );
      defparam ii1552.CONFIG_DATA = 16'h5555;
      defparam ii1552.PLACE_LOCATION = "NONE";
      defparam ii1552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1553 ( .DX(nn1553), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_649_), .F2(dummy_abc_650_), .F3(dummy_abc_651_) );
      defparam ii1553.CONFIG_DATA = 16'h5555;
      defparam ii1553.PLACE_LOCATION = "NONE";
      defparam ii1553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1554 ( .DX(nn1554), .F0(dummy_abc_652_), .F1(dummy_abc_653_), .F2(dummy_abc_654_), .F3(dummy_abc_655_) );
      defparam ii1554.CONFIG_DATA = 16'hFFFF;
      defparam ii1554.PLACE_LOCATION = "NONE";
      defparam ii1554.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_261_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_546_ ), 
        .DX( {nn1554, nn1553, nn1552, nn1551, nn1550, nn1549, nn1548, nn1547, 
              nn1546, nn1545, nn1544, nn1543, nn1542, nn1541, nn1540, nn1539, 
              nn1538, nn1537} ), 
        .SUM( {\coefcal1_divide_inst2_u120_XORCI_17|SUM_net , dummy_547_, 
              dummy_548_, dummy_549_, dummy_550_, dummy_551_, dummy_552_, dummy_553_, 
              dummy_554_, dummy_555_, dummy_556_, dummy_557_, dummy_558_, dummy_559_, 
              dummy_560_, dummy_561_, dummy_562_, dummy_563_} )
      );
    CS_LUT4_PRIM ii1575 ( .DX(nn1575), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_656_), .F3(dummy_abc_657_) );
      defparam ii1575.CONFIG_DATA = 16'h9999;
      defparam ii1575.PLACE_LOCATION = "NONE";
      defparam ii1575.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1576 ( .DX(nn1576), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[1]|Q_net ), .F2(dummy_abc_658_), .F3(dummy_abc_659_) );
      defparam ii1576.CONFIG_DATA = 16'h9999;
      defparam ii1576.PLACE_LOCATION = "NONE";
      defparam ii1576.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1577 ( .DX(nn1577), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_abc_660_), .F2(dummy_abc_661_), .F3(dummy_abc_662_) );
      defparam ii1577.CONFIG_DATA = 16'h5555;
      defparam ii1577.PLACE_LOCATION = "NONE";
      defparam ii1577.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1578 ( .DX(nn1578), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_663_), .F2(dummy_abc_664_), .F3(dummy_abc_665_) );
      defparam ii1578.CONFIG_DATA = 16'h5555;
      defparam ii1578.PLACE_LOCATION = "NONE";
      defparam ii1578.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1579 ( .DX(nn1579), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_666_), .F2(dummy_abc_667_), .F3(dummy_abc_668_) );
      defparam ii1579.CONFIG_DATA = 16'h5555;
      defparam ii1579.PLACE_LOCATION = "NONE";
      defparam ii1579.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1580 ( .DX(nn1580), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_669_), .F2(dummy_abc_670_), .F3(dummy_abc_671_) );
      defparam ii1580.CONFIG_DATA = 16'h5555;
      defparam ii1580.PLACE_LOCATION = "NONE";
      defparam ii1580.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1581 ( .DX(nn1581), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_672_), .F2(dummy_abc_673_), .F3(dummy_abc_674_) );
      defparam ii1581.CONFIG_DATA = 16'h5555;
      defparam ii1581.PLACE_LOCATION = "NONE";
      defparam ii1581.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1582 ( .DX(nn1582), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_675_), .F2(dummy_abc_676_), .F3(dummy_abc_677_) );
      defparam ii1582.CONFIG_DATA = 16'h5555;
      defparam ii1582.PLACE_LOCATION = "NONE";
      defparam ii1582.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1583 ( .DX(nn1583), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_678_), .F2(dummy_abc_679_), .F3(dummy_abc_680_) );
      defparam ii1583.CONFIG_DATA = 16'h5555;
      defparam ii1583.PLACE_LOCATION = "NONE";
      defparam ii1583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1584 ( .DX(nn1584), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_681_), .F2(dummy_abc_682_), .F3(dummy_abc_683_) );
      defparam ii1584.CONFIG_DATA = 16'h5555;
      defparam ii1584.PLACE_LOCATION = "NONE";
      defparam ii1584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1585 ( .DX(nn1585), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_684_), .F2(dummy_abc_685_), .F3(dummy_abc_686_) );
      defparam ii1585.CONFIG_DATA = 16'h5555;
      defparam ii1585.PLACE_LOCATION = "NONE";
      defparam ii1585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1586 ( .DX(nn1586), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_687_), .F2(dummy_abc_688_), .F3(dummy_abc_689_) );
      defparam ii1586.CONFIG_DATA = 16'h5555;
      defparam ii1586.PLACE_LOCATION = "NONE";
      defparam ii1586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1587 ( .DX(nn1587), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_690_), .F2(dummy_abc_691_), .F3(dummy_abc_692_) );
      defparam ii1587.CONFIG_DATA = 16'h5555;
      defparam ii1587.PLACE_LOCATION = "NONE";
      defparam ii1587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1588 ( .DX(nn1588), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_693_), .F2(dummy_abc_694_), .F3(dummy_abc_695_) );
      defparam ii1588.CONFIG_DATA = 16'h5555;
      defparam ii1588.PLACE_LOCATION = "NONE";
      defparam ii1588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1589 ( .DX(nn1589), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_696_), .F2(dummy_abc_697_), .F3(dummy_abc_698_) );
      defparam ii1589.CONFIG_DATA = 16'h5555;
      defparam ii1589.PLACE_LOCATION = "NONE";
      defparam ii1589.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1590 ( .DX(nn1590), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_699_), .F2(dummy_abc_700_), .F3(dummy_abc_701_) );
      defparam ii1590.CONFIG_DATA = 16'h5555;
      defparam ii1590.PLACE_LOCATION = "NONE";
      defparam ii1590.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1591 ( .DX(nn1591), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_702_), .F2(dummy_abc_703_), .F3(dummy_abc_704_) );
      defparam ii1591.CONFIG_DATA = 16'h5555;
      defparam ii1591.PLACE_LOCATION = "NONE";
      defparam ii1591.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_245_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, \coefcal1_yDividend__reg[16]|Q_net , 
              \coefcal1_yDividend__reg[15]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_171_ ), 
        .DX( {nn1591, nn1590, nn1589, nn1588, nn1587, nn1586, nn1585, nn1584, 
              nn1583, nn1582, nn1581, nn1580, nn1579, nn1578, nn1577, nn1576, 
              nn1575} ), 
        .SUM( {dummy_172_, \coefcal1_divide_inst2_u102_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_14|SUM_net , \coefcal1_divide_inst2_u102_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_12|SUM_net , \coefcal1_divide_inst2_u102_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_10|SUM_net , \coefcal1_divide_inst2_u102_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_8|SUM_net , \coefcal1_divide_inst2_u102_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_6|SUM_net , \coefcal1_divide_inst2_u102_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_4|SUM_net , \coefcal1_divide_inst2_u102_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_2|SUM_net , \coefcal1_divide_inst2_u102_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u102_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1611 ( .DX(nn1611), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(dummy_546_), .F2(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ), .F3(dummy_abc_705_) );
      defparam ii1611.CONFIG_DATA = 16'hB8B8;
      defparam ii1611.PLACE_LOCATION = "NONE";
      defparam ii1611.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1612 ( .DX(nn1612), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_706_), .F3(dummy_abc_707_) );
      defparam ii1612.CONFIG_DATA = 16'h9999;
      defparam ii1612.PLACE_LOCATION = "NONE";
      defparam ii1612.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1613 ( .DX(nn1613), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_546_) );
      defparam ii1613.CONFIG_DATA = 16'hA569;
      defparam ii1613.PLACE_LOCATION = "NONE";
      defparam ii1613.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1614 ( .DX(nn1614), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_546_), .F3(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ) );
      defparam ii1614.CONFIG_DATA = 16'h9C93;
      defparam ii1614.PLACE_LOCATION = "NONE";
      defparam ii1614.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1615 ( .DX(nn1615), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_708_), .F2(dummy_abc_709_), .F3(dummy_abc_710_) );
      defparam ii1615.CONFIG_DATA = 16'h5555;
      defparam ii1615.PLACE_LOCATION = "NONE";
      defparam ii1615.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1616 ( .DX(nn1616), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_711_), .F2(dummy_abc_712_), .F3(dummy_abc_713_) );
      defparam ii1616.CONFIG_DATA = 16'h5555;
      defparam ii1616.PLACE_LOCATION = "NONE";
      defparam ii1616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1617 ( .DX(nn1617), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_714_), .F2(dummy_abc_715_), .F3(dummy_abc_716_) );
      defparam ii1617.CONFIG_DATA = 16'h5555;
      defparam ii1617.PLACE_LOCATION = "NONE";
      defparam ii1617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1618 ( .DX(nn1618), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_717_), .F2(dummy_abc_718_), .F3(dummy_abc_719_) );
      defparam ii1618.CONFIG_DATA = 16'h5555;
      defparam ii1618.PLACE_LOCATION = "NONE";
      defparam ii1618.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1619 ( .DX(nn1619), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_720_), .F2(dummy_abc_721_), .F3(dummy_abc_722_) );
      defparam ii1619.CONFIG_DATA = 16'h5555;
      defparam ii1619.PLACE_LOCATION = "NONE";
      defparam ii1619.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1620 ( .DX(nn1620), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_723_), .F2(dummy_abc_724_), .F3(dummy_abc_725_) );
      defparam ii1620.CONFIG_DATA = 16'h5555;
      defparam ii1620.PLACE_LOCATION = "NONE";
      defparam ii1620.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1621 ( .DX(nn1621), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_726_), .F2(dummy_abc_727_), .F3(dummy_abc_728_) );
      defparam ii1621.CONFIG_DATA = 16'h5555;
      defparam ii1621.PLACE_LOCATION = "NONE";
      defparam ii1621.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1622 ( .DX(nn1622), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_729_), .F2(dummy_abc_730_), .F3(dummy_abc_731_) );
      defparam ii1622.CONFIG_DATA = 16'h5555;
      defparam ii1622.PLACE_LOCATION = "NONE";
      defparam ii1622.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1623 ( .DX(nn1623), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_732_), .F2(dummy_abc_733_), .F3(dummy_abc_734_) );
      defparam ii1623.CONFIG_DATA = 16'h5555;
      defparam ii1623.PLACE_LOCATION = "NONE";
      defparam ii1623.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1624 ( .DX(nn1624), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_735_), .F2(dummy_abc_736_), .F3(dummy_abc_737_) );
      defparam ii1624.CONFIG_DATA = 16'h5555;
      defparam ii1624.PLACE_LOCATION = "NONE";
      defparam ii1624.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1625 ( .DX(nn1625), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_738_), .F2(dummy_abc_739_), .F3(dummy_abc_740_) );
      defparam ii1625.CONFIG_DATA = 16'h5555;
      defparam ii1625.PLACE_LOCATION = "NONE";
      defparam ii1625.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1626 ( .DX(nn1626), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_741_), .F2(dummy_abc_742_), .F3(dummy_abc_743_) );
      defparam ii1626.CONFIG_DATA = 16'h5555;
      defparam ii1626.PLACE_LOCATION = "NONE";
      defparam ii1626.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1627 ( .DX(nn1627), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_744_), .F2(dummy_abc_745_), .F3(dummy_abc_746_) );
      defparam ii1627.CONFIG_DATA = 16'h5555;
      defparam ii1627.PLACE_LOCATION = "NONE";
      defparam ii1627.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1628 ( .DX(nn1628), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_747_), .F2(dummy_abc_748_), .F3(dummy_abc_749_) );
      defparam ii1628.CONFIG_DATA = 16'h5555;
      defparam ii1628.PLACE_LOCATION = "NONE";
      defparam ii1628.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1629 ( .DX(nn1629), .F0(dummy_abc_750_), .F1(dummy_abc_751_), .F2(dummy_abc_752_), .F3(dummy_abc_753_) );
      defparam ii1629.CONFIG_DATA = 16'hFFFF;
      defparam ii1629.PLACE_LOCATION = "NONE";
      defparam ii1629.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_262_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_565_ ), 
        .DX( {nn1629, nn1628, nn1627, nn1626, nn1625, nn1624, nn1623, nn1622, 
              nn1621, nn1620, nn1619, nn1618, nn1617, nn1616, nn1615, nn1614, 
              nn1613, nn1612} ), 
        .SUM( {\coefcal1_divide_inst2_u122_XORCI_17|SUM_net , dummy_566_, 
              dummy_567_, dummy_568_, dummy_569_, dummy_570_, dummy_571_, dummy_572_, 
              dummy_573_, dummy_574_, dummy_575_, dummy_576_, dummy_577_, dummy_578_, 
              dummy_579_, dummy_580_, dummy_581_, dummy_582_} )
      );
    CS_LUT4_PRIM ii1650 ( .DX(nn1650), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_546_), .F3(dummy_abc_754_) );
      defparam ii1650.CONFIG_DATA = 16'hA6A6;
      defparam ii1650.PLACE_LOCATION = "NONE";
      defparam ii1650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1651 ( .DX(nn1651), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_755_), .F3(dummy_abc_756_) );
      defparam ii1651.CONFIG_DATA = 16'h9999;
      defparam ii1651.PLACE_LOCATION = "NONE";
      defparam ii1651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1652 ( .DX(nn1652), .F0(\coefcal1_yDividend__reg[15]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_546_) );
      defparam ii1652.CONFIG_DATA = 16'hA569;
      defparam ii1652.PLACE_LOCATION = "NONE";
      defparam ii1652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1653 ( .DX(nn1653), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(dummy_546_), .F3(\coefcal1_divide_inst2_u102_XORCI_1|SUM_net ) );
      defparam ii1653.CONFIG_DATA = 16'h9C93;
      defparam ii1653.PLACE_LOCATION = "NONE";
      defparam ii1653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1654 ( .DX(nn1654), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(dummy_abc_757_), .F2(dummy_abc_758_), .F3(dummy_abc_759_) );
      defparam ii1654.CONFIG_DATA = 16'h5555;
      defparam ii1654.PLACE_LOCATION = "NONE";
      defparam ii1654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1655 ( .DX(nn1655), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_760_), .F2(dummy_abc_761_), .F3(dummy_abc_762_) );
      defparam ii1655.CONFIG_DATA = 16'h5555;
      defparam ii1655.PLACE_LOCATION = "NONE";
      defparam ii1655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1656 ( .DX(nn1656), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_763_), .F2(dummy_abc_764_), .F3(dummy_abc_765_) );
      defparam ii1656.CONFIG_DATA = 16'h5555;
      defparam ii1656.PLACE_LOCATION = "NONE";
      defparam ii1656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1657 ( .DX(nn1657), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_766_), .F2(dummy_abc_767_), .F3(dummy_abc_768_) );
      defparam ii1657.CONFIG_DATA = 16'h5555;
      defparam ii1657.PLACE_LOCATION = "NONE";
      defparam ii1657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1658 ( .DX(nn1658), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_769_), .F2(dummy_abc_770_), .F3(dummy_abc_771_) );
      defparam ii1658.CONFIG_DATA = 16'h5555;
      defparam ii1658.PLACE_LOCATION = "NONE";
      defparam ii1658.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1659 ( .DX(nn1659), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_772_), .F2(dummy_abc_773_), .F3(dummy_abc_774_) );
      defparam ii1659.CONFIG_DATA = 16'h5555;
      defparam ii1659.PLACE_LOCATION = "NONE";
      defparam ii1659.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1660 ( .DX(nn1660), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_775_), .F2(dummy_abc_776_), .F3(dummy_abc_777_) );
      defparam ii1660.CONFIG_DATA = 16'h5555;
      defparam ii1660.PLACE_LOCATION = "NONE";
      defparam ii1660.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1661 ( .DX(nn1661), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_778_), .F2(dummy_abc_779_), .F3(dummy_abc_780_) );
      defparam ii1661.CONFIG_DATA = 16'h5555;
      defparam ii1661.PLACE_LOCATION = "NONE";
      defparam ii1661.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1662 ( .DX(nn1662), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_781_), .F2(dummy_abc_782_), .F3(dummy_abc_783_) );
      defparam ii1662.CONFIG_DATA = 16'h5555;
      defparam ii1662.PLACE_LOCATION = "NONE";
      defparam ii1662.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1663 ( .DX(nn1663), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_784_), .F2(dummy_abc_785_), .F3(dummy_abc_786_) );
      defparam ii1663.CONFIG_DATA = 16'h5555;
      defparam ii1663.PLACE_LOCATION = "NONE";
      defparam ii1663.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1664 ( .DX(nn1664), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_787_), .F2(dummy_abc_788_), .F3(dummy_abc_789_) );
      defparam ii1664.CONFIG_DATA = 16'h5555;
      defparam ii1664.PLACE_LOCATION = "NONE";
      defparam ii1664.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1665 ( .DX(nn1665), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_790_), .F2(dummy_abc_791_), .F3(dummy_abc_792_) );
      defparam ii1665.CONFIG_DATA = 16'h5555;
      defparam ii1665.PLACE_LOCATION = "NONE";
      defparam ii1665.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1666 ( .DX(nn1666), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_793_), .F2(dummy_abc_794_), .F3(dummy_abc_795_) );
      defparam ii1666.CONFIG_DATA = 16'h5555;
      defparam ii1666.PLACE_LOCATION = "NONE";
      defparam ii1666.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1667 ( .DX(nn1667), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_796_), .F2(dummy_abc_797_), .F3(dummy_abc_798_) );
      defparam ii1667.CONFIG_DATA = 16'h5555;
      defparam ii1667.PLACE_LOCATION = "NONE";
      defparam ii1667.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_246_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn1611, 
              nn1650, \coefcal1_yDividend__reg[14]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_173_ ), 
        .DX( {nn1667, nn1666, nn1665, nn1664, nn1663, nn1662, nn1661, nn1660, 
              nn1659, nn1658, nn1657, nn1656, nn1655, nn1654, nn1653, nn1652, 
              nn1651} ), 
        .SUM( {dummy_174_, \coefcal1_divide_inst2_u103_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_14|SUM_net , \coefcal1_divide_inst2_u103_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_12|SUM_net , \coefcal1_divide_inst2_u103_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_10|SUM_net , \coefcal1_divide_inst2_u103_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_8|SUM_net , \coefcal1_divide_inst2_u103_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_6|SUM_net , \coefcal1_divide_inst2_u103_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_4|SUM_net , \coefcal1_divide_inst2_u103_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_2|SUM_net , \coefcal1_divide_inst2_u103_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u103_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1687 ( .DX(nn1687), .F0(nn1611), .F1(dummy_565_), .F2(\coefcal1_divide_inst2_u103_XORCI_2|SUM_net ), .F3(dummy_abc_799_) );
      defparam ii1687.CONFIG_DATA = 16'hB8B8;
      defparam ii1687.PLACE_LOCATION = "NONE";
      defparam ii1687.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1688 ( .DX(nn1688), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_800_), .F3(dummy_abc_801_) );
      defparam ii1688.CONFIG_DATA = 16'h9999;
      defparam ii1688.PLACE_LOCATION = "NONE";
      defparam ii1688.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1689 ( .DX(nn1689), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_565_) );
      defparam ii1689.CONFIG_DATA = 16'hA569;
      defparam ii1689.PLACE_LOCATION = "NONE";
      defparam ii1689.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1690 ( .DX(nn1690), .F0(dummy_565_), .F1(nn1650), .F2(\coefcal1_divide_inst2_u103_XORCI_1|SUM_net ), .F3(dummy_abc_802_) );
      defparam ii1690.CONFIG_DATA = 16'hD8D8;
      defparam ii1690.PLACE_LOCATION = "NONE";
      defparam ii1690.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1691 ( .DX(nn1691), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1690), .F2(dummy_abc_803_), .F3(dummy_abc_804_) );
      defparam ii1691.CONFIG_DATA = 16'h9999;
      defparam ii1691.PLACE_LOCATION = "NONE";
      defparam ii1691.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1692 ( .DX(nn1692), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1687), .F2(dummy_abc_805_), .F3(dummy_abc_806_) );
      defparam ii1692.CONFIG_DATA = 16'h9999;
      defparam ii1692.PLACE_LOCATION = "NONE";
      defparam ii1692.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1693 ( .DX(nn1693), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_807_), .F2(dummy_abc_808_), .F3(dummy_abc_809_) );
      defparam ii1693.CONFIG_DATA = 16'h5555;
      defparam ii1693.PLACE_LOCATION = "NONE";
      defparam ii1693.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1694 ( .DX(nn1694), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_810_), .F2(dummy_abc_811_), .F3(dummy_abc_812_) );
      defparam ii1694.CONFIG_DATA = 16'h5555;
      defparam ii1694.PLACE_LOCATION = "NONE";
      defparam ii1694.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1695 ( .DX(nn1695), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_813_), .F2(dummy_abc_814_), .F3(dummy_abc_815_) );
      defparam ii1695.CONFIG_DATA = 16'h5555;
      defparam ii1695.PLACE_LOCATION = "NONE";
      defparam ii1695.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1696 ( .DX(nn1696), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_816_), .F2(dummy_abc_817_), .F3(dummy_abc_818_) );
      defparam ii1696.CONFIG_DATA = 16'h5555;
      defparam ii1696.PLACE_LOCATION = "NONE";
      defparam ii1696.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1697 ( .DX(nn1697), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_819_), .F2(dummy_abc_820_), .F3(dummy_abc_821_) );
      defparam ii1697.CONFIG_DATA = 16'h5555;
      defparam ii1697.PLACE_LOCATION = "NONE";
      defparam ii1697.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1698 ( .DX(nn1698), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_822_), .F2(dummy_abc_823_), .F3(dummy_abc_824_) );
      defparam ii1698.CONFIG_DATA = 16'h5555;
      defparam ii1698.PLACE_LOCATION = "NONE";
      defparam ii1698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1699 ( .DX(nn1699), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_825_), .F2(dummy_abc_826_), .F3(dummy_abc_827_) );
      defparam ii1699.CONFIG_DATA = 16'h5555;
      defparam ii1699.PLACE_LOCATION = "NONE";
      defparam ii1699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1700 ( .DX(nn1700), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_828_), .F2(dummy_abc_829_), .F3(dummy_abc_830_) );
      defparam ii1700.CONFIG_DATA = 16'h5555;
      defparam ii1700.PLACE_LOCATION = "NONE";
      defparam ii1700.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1701 ( .DX(nn1701), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_831_), .F2(dummy_abc_832_), .F3(dummy_abc_833_) );
      defparam ii1701.CONFIG_DATA = 16'h5555;
      defparam ii1701.PLACE_LOCATION = "NONE";
      defparam ii1701.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1702 ( .DX(nn1702), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_834_), .F2(dummy_abc_835_), .F3(dummy_abc_836_) );
      defparam ii1702.CONFIG_DATA = 16'h5555;
      defparam ii1702.PLACE_LOCATION = "NONE";
      defparam ii1702.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1703 ( .DX(nn1703), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_837_), .F2(dummy_abc_838_), .F3(dummy_abc_839_) );
      defparam ii1703.CONFIG_DATA = 16'h5555;
      defparam ii1703.PLACE_LOCATION = "NONE";
      defparam ii1703.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1704 ( .DX(nn1704), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_840_), .F2(dummy_abc_841_), .F3(dummy_abc_842_) );
      defparam ii1704.CONFIG_DATA = 16'h5555;
      defparam ii1704.PLACE_LOCATION = "NONE";
      defparam ii1704.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1705 ( .DX(nn1705), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_843_), .F2(dummy_abc_844_), .F3(dummy_abc_845_) );
      defparam ii1705.CONFIG_DATA = 16'h5555;
      defparam ii1705.PLACE_LOCATION = "NONE";
      defparam ii1705.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1706 ( .DX(nn1706), .F0(dummy_abc_846_), .F1(dummy_abc_847_), .F2(dummy_abc_848_), .F3(dummy_abc_849_) );
      defparam ii1706.CONFIG_DATA = 16'hFFFF;
      defparam ii1706.PLACE_LOCATION = "NONE";
      defparam ii1706.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_263_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_584_ ), 
        .DX( {nn1706, nn1705, nn1704, nn1703, nn1702, nn1701, nn1700, nn1699, 
              nn1698, nn1697, nn1696, nn1695, nn1694, nn1693, nn1692, nn1691, 
              nn1689, nn1688} ), 
        .SUM( {\coefcal1_divide_inst2_u124_XORCI_17|SUM_net , dummy_585_, 
              dummy_586_, dummy_587_, dummy_588_, dummy_589_, dummy_590_, dummy_591_, 
              dummy_592_, dummy_593_, dummy_594_, dummy_595_, dummy_596_, dummy_597_, 
              dummy_598_, dummy_599_, dummy_600_, dummy_601_} )
      );
    CS_LUT4_PRIM ii1727 ( .DX(nn1727), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_565_), .F3(dummy_abc_850_) );
      defparam ii1727.CONFIG_DATA = 16'hA6A6;
      defparam ii1727.PLACE_LOCATION = "NONE";
      defparam ii1727.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1728 ( .DX(nn1728), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_851_), .F3(dummy_abc_852_) );
      defparam ii1728.CONFIG_DATA = 16'h9999;
      defparam ii1728.PLACE_LOCATION = "NONE";
      defparam ii1728.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1729 ( .DX(nn1729), .F0(\coefcal1_yDividend__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_565_) );
      defparam ii1729.CONFIG_DATA = 16'hA569;
      defparam ii1729.PLACE_LOCATION = "NONE";
      defparam ii1729.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1730 ( .DX(nn1730), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1690), .F2(dummy_abc_853_), .F3(dummy_abc_854_) );
      defparam ii1730.CONFIG_DATA = 16'h9999;
      defparam ii1730.PLACE_LOCATION = "NONE";
      defparam ii1730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1731 ( .DX(nn1731), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1687), .F2(dummy_abc_855_), .F3(dummy_abc_856_) );
      defparam ii1731.CONFIG_DATA = 16'h9999;
      defparam ii1731.PLACE_LOCATION = "NONE";
      defparam ii1731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1732 ( .DX(nn1732), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(dummy_abc_857_), .F2(dummy_abc_858_), .F3(dummy_abc_859_) );
      defparam ii1732.CONFIG_DATA = 16'h5555;
      defparam ii1732.PLACE_LOCATION = "NONE";
      defparam ii1732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1733 ( .DX(nn1733), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_860_), .F2(dummy_abc_861_), .F3(dummy_abc_862_) );
      defparam ii1733.CONFIG_DATA = 16'h5555;
      defparam ii1733.PLACE_LOCATION = "NONE";
      defparam ii1733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1734 ( .DX(nn1734), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_863_), .F2(dummy_abc_864_), .F3(dummy_abc_865_) );
      defparam ii1734.CONFIG_DATA = 16'h5555;
      defparam ii1734.PLACE_LOCATION = "NONE";
      defparam ii1734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1735 ( .DX(nn1735), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_866_), .F2(dummy_abc_867_), .F3(dummy_abc_868_) );
      defparam ii1735.CONFIG_DATA = 16'h5555;
      defparam ii1735.PLACE_LOCATION = "NONE";
      defparam ii1735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1736 ( .DX(nn1736), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_869_), .F2(dummy_abc_870_), .F3(dummy_abc_871_) );
      defparam ii1736.CONFIG_DATA = 16'h5555;
      defparam ii1736.PLACE_LOCATION = "NONE";
      defparam ii1736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1737 ( .DX(nn1737), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_872_), .F2(dummy_abc_873_), .F3(dummy_abc_874_) );
      defparam ii1737.CONFIG_DATA = 16'h5555;
      defparam ii1737.PLACE_LOCATION = "NONE";
      defparam ii1737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1738 ( .DX(nn1738), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_875_), .F2(dummy_abc_876_), .F3(dummy_abc_877_) );
      defparam ii1738.CONFIG_DATA = 16'h5555;
      defparam ii1738.PLACE_LOCATION = "NONE";
      defparam ii1738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1739 ( .DX(nn1739), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_878_), .F2(dummy_abc_879_), .F3(dummy_abc_880_) );
      defparam ii1739.CONFIG_DATA = 16'h5555;
      defparam ii1739.PLACE_LOCATION = "NONE";
      defparam ii1739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1740 ( .DX(nn1740), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_881_), .F2(dummy_abc_882_), .F3(dummy_abc_883_) );
      defparam ii1740.CONFIG_DATA = 16'h5555;
      defparam ii1740.PLACE_LOCATION = "NONE";
      defparam ii1740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1741 ( .DX(nn1741), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_884_), .F2(dummy_abc_885_), .F3(dummy_abc_886_) );
      defparam ii1741.CONFIG_DATA = 16'h5555;
      defparam ii1741.PLACE_LOCATION = "NONE";
      defparam ii1741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1742 ( .DX(nn1742), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_887_), .F2(dummy_abc_888_), .F3(dummy_abc_889_) );
      defparam ii1742.CONFIG_DATA = 16'h5555;
      defparam ii1742.PLACE_LOCATION = "NONE";
      defparam ii1742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1743 ( .DX(nn1743), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_890_), .F2(dummy_abc_891_), .F3(dummy_abc_892_) );
      defparam ii1743.CONFIG_DATA = 16'h5555;
      defparam ii1743.PLACE_LOCATION = "NONE";
      defparam ii1743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1744 ( .DX(nn1744), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_893_), .F2(dummy_abc_894_), .F3(dummy_abc_895_) );
      defparam ii1744.CONFIG_DATA = 16'h5555;
      defparam ii1744.PLACE_LOCATION = "NONE";
      defparam ii1744.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_247_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn1687, nn1690, nn1727, 
              \coefcal1_yDividend__reg[13]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_175_ ), 
        .DX( {nn1744, nn1743, nn1742, nn1741, nn1740, nn1739, nn1738, nn1737, 
              nn1736, nn1735, nn1734, nn1733, nn1732, nn1731, nn1730, nn1729, 
              nn1728} ), 
        .SUM( {dummy_176_, \coefcal1_divide_inst2_u104_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_14|SUM_net , \coefcal1_divide_inst2_u104_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_12|SUM_net , \coefcal1_divide_inst2_u104_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_10|SUM_net , \coefcal1_divide_inst2_u104_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_8|SUM_net , \coefcal1_divide_inst2_u104_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_6|SUM_net , \coefcal1_divide_inst2_u104_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_4|SUM_net , \coefcal1_divide_inst2_u104_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_2|SUM_net , \coefcal1_divide_inst2_u104_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u104_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1764 ( .DX(nn1764), .F0(nn1687), .F1(dummy_584_), .F2(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ), .F3(dummy_abc_896_) );
      defparam ii1764.CONFIG_DATA = 16'hB8B8;
      defparam ii1764.PLACE_LOCATION = "NONE";
      defparam ii1764.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1765 ( .DX(nn1765), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_897_), .F3(dummy_abc_898_) );
      defparam ii1765.CONFIG_DATA = 16'h9999;
      defparam ii1765.PLACE_LOCATION = "NONE";
      defparam ii1765.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1766 ( .DX(nn1766), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_584_) );
      defparam ii1766.CONFIG_DATA = 16'hA569;
      defparam ii1766.PLACE_LOCATION = "NONE";
      defparam ii1766.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1767 ( .DX(nn1767), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_584_), .F2(nn1727), .F3(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ) );
      defparam ii1767.CONFIG_DATA = 16'hA695;
      defparam ii1767.PLACE_LOCATION = "NONE";
      defparam ii1767.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1768 ( .DX(nn1768), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1690), .F2(dummy_584_), .F3(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ) );
      defparam ii1768.CONFIG_DATA = 16'h9A95;
      defparam ii1768.PLACE_LOCATION = "NONE";
      defparam ii1768.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1769 ( .DX(nn1769), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1687), .F2(dummy_584_), .F3(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ) );
      defparam ii1769.CONFIG_DATA = 16'h9A95;
      defparam ii1769.PLACE_LOCATION = "NONE";
      defparam ii1769.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1770 ( .DX(nn1770), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_899_), .F2(dummy_abc_900_), .F3(dummy_abc_901_) );
      defparam ii1770.CONFIG_DATA = 16'h5555;
      defparam ii1770.PLACE_LOCATION = "NONE";
      defparam ii1770.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1771 ( .DX(nn1771), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_902_), .F2(dummy_abc_903_), .F3(dummy_abc_904_) );
      defparam ii1771.CONFIG_DATA = 16'h5555;
      defparam ii1771.PLACE_LOCATION = "NONE";
      defparam ii1771.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1772 ( .DX(nn1772), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_905_), .F2(dummy_abc_906_), .F3(dummy_abc_907_) );
      defparam ii1772.CONFIG_DATA = 16'h5555;
      defparam ii1772.PLACE_LOCATION = "NONE";
      defparam ii1772.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1773 ( .DX(nn1773), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_908_), .F2(dummy_abc_909_), .F3(dummy_abc_910_) );
      defparam ii1773.CONFIG_DATA = 16'h5555;
      defparam ii1773.PLACE_LOCATION = "NONE";
      defparam ii1773.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1774 ( .DX(nn1774), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_911_), .F2(dummy_abc_912_), .F3(dummy_abc_913_) );
      defparam ii1774.CONFIG_DATA = 16'h5555;
      defparam ii1774.PLACE_LOCATION = "NONE";
      defparam ii1774.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1775 ( .DX(nn1775), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_914_), .F2(dummy_abc_915_), .F3(dummy_abc_916_) );
      defparam ii1775.CONFIG_DATA = 16'h5555;
      defparam ii1775.PLACE_LOCATION = "NONE";
      defparam ii1775.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1776 ( .DX(nn1776), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_917_), .F2(dummy_abc_918_), .F3(dummy_abc_919_) );
      defparam ii1776.CONFIG_DATA = 16'h5555;
      defparam ii1776.PLACE_LOCATION = "NONE";
      defparam ii1776.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1777 ( .DX(nn1777), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_920_), .F2(dummy_abc_921_), .F3(dummy_abc_922_) );
      defparam ii1777.CONFIG_DATA = 16'h5555;
      defparam ii1777.PLACE_LOCATION = "NONE";
      defparam ii1777.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1778 ( .DX(nn1778), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_923_), .F2(dummy_abc_924_), .F3(dummy_abc_925_) );
      defparam ii1778.CONFIG_DATA = 16'h5555;
      defparam ii1778.PLACE_LOCATION = "NONE";
      defparam ii1778.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1779 ( .DX(nn1779), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_926_), .F2(dummy_abc_927_), .F3(dummy_abc_928_) );
      defparam ii1779.CONFIG_DATA = 16'h5555;
      defparam ii1779.PLACE_LOCATION = "NONE";
      defparam ii1779.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1780 ( .DX(nn1780), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_929_), .F2(dummy_abc_930_), .F3(dummy_abc_931_) );
      defparam ii1780.CONFIG_DATA = 16'h5555;
      defparam ii1780.PLACE_LOCATION = "NONE";
      defparam ii1780.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1781 ( .DX(nn1781), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_932_), .F2(dummy_abc_933_), .F3(dummy_abc_934_) );
      defparam ii1781.CONFIG_DATA = 16'h5555;
      defparam ii1781.PLACE_LOCATION = "NONE";
      defparam ii1781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1782 ( .DX(nn1782), .F0(dummy_abc_935_), .F1(dummy_abc_936_), .F2(dummy_abc_937_), .F3(dummy_abc_938_) );
      defparam ii1782.CONFIG_DATA = 16'hFFFF;
      defparam ii1782.PLACE_LOCATION = "NONE";
      defparam ii1782.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_264_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_603_ ), 
        .DX( {nn1782, nn1781, nn1780, nn1779, nn1778, nn1777, nn1776, nn1775, 
              nn1774, nn1773, nn1772, nn1771, nn1770, nn1769, nn1768, nn1767, 
              nn1766, nn1765} ), 
        .SUM( {\coefcal1_divide_inst2_u126_XORCI_17|SUM_net , dummy_604_, 
              dummy_605_, dummy_606_, dummy_607_, dummy_608_, dummy_609_, dummy_610_, 
              dummy_611_, dummy_612_, dummy_613_, dummy_614_, dummy_615_, dummy_616_, 
              dummy_617_, dummy_618_, dummy_619_, dummy_620_} )
      );
    CS_LUT4_PRIM ii1803 ( .DX(nn1803), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_584_), .F3(dummy_abc_939_) );
      defparam ii1803.CONFIG_DATA = 16'hA6A6;
      defparam ii1803.PLACE_LOCATION = "NONE";
      defparam ii1803.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1804 ( .DX(nn1804), .F0(dummy_584_), .F1(nn1727), .F2(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ), .F3(dummy_abc_940_) );
      defparam ii1804.CONFIG_DATA = 16'hD8D8;
      defparam ii1804.PLACE_LOCATION = "NONE";
      defparam ii1804.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1805 ( .DX(nn1805), .F0(nn1690), .F1(dummy_584_), .F2(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ), .F3(dummy_abc_941_) );
      defparam ii1805.CONFIG_DATA = 16'hB8B8;
      defparam ii1805.PLACE_LOCATION = "NONE";
      defparam ii1805.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1806 ( .DX(nn1806), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_942_), .F3(dummy_abc_943_) );
      defparam ii1806.CONFIG_DATA = 16'h9999;
      defparam ii1806.PLACE_LOCATION = "NONE";
      defparam ii1806.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1807 ( .DX(nn1807), .F0(\coefcal1_yDividend__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_584_) );
      defparam ii1807.CONFIG_DATA = 16'hA569;
      defparam ii1807.PLACE_LOCATION = "NONE";
      defparam ii1807.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1808 ( .DX(nn1808), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_584_), .F2(nn1727), .F3(\coefcal1_divide_inst2_u104_XORCI_1|SUM_net ) );
      defparam ii1808.CONFIG_DATA = 16'hA695;
      defparam ii1808.PLACE_LOCATION = "NONE";
      defparam ii1808.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1809 ( .DX(nn1809), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1690), .F2(dummy_584_), .F3(\coefcal1_divide_inst2_u104_XORCI_2|SUM_net ) );
      defparam ii1809.CONFIG_DATA = 16'h9A95;
      defparam ii1809.PLACE_LOCATION = "NONE";
      defparam ii1809.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1810 ( .DX(nn1810), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1687), .F2(dummy_584_), .F3(\coefcal1_divide_inst2_u104_XORCI_3|SUM_net ) );
      defparam ii1810.CONFIG_DATA = 16'h9A95;
      defparam ii1810.PLACE_LOCATION = "NONE";
      defparam ii1810.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1811 ( .DX(nn1811), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(dummy_abc_944_), .F2(dummy_abc_945_), .F3(dummy_abc_946_) );
      defparam ii1811.CONFIG_DATA = 16'h5555;
      defparam ii1811.PLACE_LOCATION = "NONE";
      defparam ii1811.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1812 ( .DX(nn1812), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_947_), .F2(dummy_abc_948_), .F3(dummy_abc_949_) );
      defparam ii1812.CONFIG_DATA = 16'h5555;
      defparam ii1812.PLACE_LOCATION = "NONE";
      defparam ii1812.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1813 ( .DX(nn1813), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_950_), .F2(dummy_abc_951_), .F3(dummy_abc_952_) );
      defparam ii1813.CONFIG_DATA = 16'h5555;
      defparam ii1813.PLACE_LOCATION = "NONE";
      defparam ii1813.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1814 ( .DX(nn1814), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_953_), .F2(dummy_abc_954_), .F3(dummy_abc_955_) );
      defparam ii1814.CONFIG_DATA = 16'h5555;
      defparam ii1814.PLACE_LOCATION = "NONE";
      defparam ii1814.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1815 ( .DX(nn1815), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_956_), .F2(dummy_abc_957_), .F3(dummy_abc_958_) );
      defparam ii1815.CONFIG_DATA = 16'h5555;
      defparam ii1815.PLACE_LOCATION = "NONE";
      defparam ii1815.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1816 ( .DX(nn1816), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_959_), .F2(dummy_abc_960_), .F3(dummy_abc_961_) );
      defparam ii1816.CONFIG_DATA = 16'h5555;
      defparam ii1816.PLACE_LOCATION = "NONE";
      defparam ii1816.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1817 ( .DX(nn1817), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_962_), .F2(dummy_abc_963_), .F3(dummy_abc_964_) );
      defparam ii1817.CONFIG_DATA = 16'h5555;
      defparam ii1817.PLACE_LOCATION = "NONE";
      defparam ii1817.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1818 ( .DX(nn1818), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_965_), .F2(dummy_abc_966_), .F3(dummy_abc_967_) );
      defparam ii1818.CONFIG_DATA = 16'h5555;
      defparam ii1818.PLACE_LOCATION = "NONE";
      defparam ii1818.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1819 ( .DX(nn1819), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_968_), .F2(dummy_abc_969_), .F3(dummy_abc_970_) );
      defparam ii1819.CONFIG_DATA = 16'h5555;
      defparam ii1819.PLACE_LOCATION = "NONE";
      defparam ii1819.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1820 ( .DX(nn1820), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_971_), .F2(dummy_abc_972_), .F3(dummy_abc_973_) );
      defparam ii1820.CONFIG_DATA = 16'h5555;
      defparam ii1820.PLACE_LOCATION = "NONE";
      defparam ii1820.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1821 ( .DX(nn1821), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_974_), .F2(dummy_abc_975_), .F3(dummy_abc_976_) );
      defparam ii1821.CONFIG_DATA = 16'h5555;
      defparam ii1821.PLACE_LOCATION = "NONE";
      defparam ii1821.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1822 ( .DX(nn1822), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_977_), .F2(dummy_abc_978_), .F3(dummy_abc_979_) );
      defparam ii1822.CONFIG_DATA = 16'h5555;
      defparam ii1822.PLACE_LOCATION = "NONE";
      defparam ii1822.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_248_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn1764, nn1805, nn1804, nn1803, 
              \coefcal1_yDividend__reg[12]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_177_ ), 
        .DX( {nn1822, nn1821, nn1820, nn1819, nn1818, nn1817, nn1816, nn1815, 
              nn1814, nn1813, nn1812, nn1811, nn1810, nn1809, nn1808, nn1807, 
              nn1806} ), 
        .SUM( {dummy_178_, \coefcal1_divide_inst2_u105_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_14|SUM_net , \coefcal1_divide_inst2_u105_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_12|SUM_net , \coefcal1_divide_inst2_u105_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_10|SUM_net , \coefcal1_divide_inst2_u105_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_8|SUM_net , \coefcal1_divide_inst2_u105_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_6|SUM_net , \coefcal1_divide_inst2_u105_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_4|SUM_net , \coefcal1_divide_inst2_u105_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_2|SUM_net , \coefcal1_divide_inst2_u105_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u105_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1842 ( .DX(nn1842), .F0(dummy_603_), .F1(\coefcal1_divide_inst2_u105_XORCI_4|SUM_net ), .F2(dummy_abc_980_), .F3(dummy_abc_981_) );
      defparam ii1842.CONFIG_DATA = 16'h1111;
      defparam ii1842.PLACE_LOCATION = "NONE";
      defparam ii1842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1843 ( .DX(nn1843), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_982_), .F3(dummy_abc_983_) );
      defparam ii1843.CONFIG_DATA = 16'h9999;
      defparam ii1843.PLACE_LOCATION = "NONE";
      defparam ii1843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1844 ( .DX(nn1844), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_603_) );
      defparam ii1844.CONFIG_DATA = 16'hA569;
      defparam ii1844.PLACE_LOCATION = "NONE";
      defparam ii1844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1845 ( .DX(nn1845), .F0(dummy_603_), .F1(nn1803), .F2(\coefcal1_divide_inst2_u105_XORCI_1|SUM_net ), .F3(dummy_abc_984_) );
      defparam ii1845.CONFIG_DATA = 16'hD8D8;
      defparam ii1845.PLACE_LOCATION = "NONE";
      defparam ii1845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1846 ( .DX(nn1846), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1845), .F2(dummy_abc_985_), .F3(dummy_abc_986_) );
      defparam ii1846.CONFIG_DATA = 16'h9999;
      defparam ii1846.PLACE_LOCATION = "NONE";
      defparam ii1846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1847 ( .DX(nn1847), .F0(nn1804), .F1(dummy_603_), .F2(\coefcal1_divide_inst2_u105_XORCI_2|SUM_net ), .F3(dummy_abc_987_) );
      defparam ii1847.CONFIG_DATA = 16'hB8B8;
      defparam ii1847.PLACE_LOCATION = "NONE";
      defparam ii1847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1848 ( .DX(nn1848), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1847), .F2(dummy_abc_988_), .F3(dummy_abc_989_) );
      defparam ii1848.CONFIG_DATA = 16'h9999;
      defparam ii1848.PLACE_LOCATION = "NONE";
      defparam ii1848.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1849 ( .DX(nn1849), .F0(nn1805), .F1(dummy_603_), .F2(\coefcal1_divide_inst2_u105_XORCI_3|SUM_net ), .F3(dummy_abc_990_) );
      defparam ii1849.CONFIG_DATA = 16'hB8B8;
      defparam ii1849.PLACE_LOCATION = "NONE";
      defparam ii1849.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1850 ( .DX(nn1850), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1849), .F2(dummy_abc_991_), .F3(dummy_abc_992_) );
      defparam ii1850.CONFIG_DATA = 16'h9999;
      defparam ii1850.PLACE_LOCATION = "NONE";
      defparam ii1850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1851 ( .DX(nn1851), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1764), .F2(nn1842), .F3(dummy_abc_993_) );
      defparam ii1851.CONFIG_DATA = 16'hD9D9;
      defparam ii1851.PLACE_LOCATION = "NONE";
      defparam ii1851.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1852 ( .DX(nn1852), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_994_), .F2(dummy_abc_995_), .F3(dummy_abc_996_) );
      defparam ii1852.CONFIG_DATA = 16'h5555;
      defparam ii1852.PLACE_LOCATION = "NONE";
      defparam ii1852.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1853 ( .DX(nn1853), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_997_), .F2(dummy_abc_998_), .F3(dummy_abc_999_) );
      defparam ii1853.CONFIG_DATA = 16'h5555;
      defparam ii1853.PLACE_LOCATION = "NONE";
      defparam ii1853.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1854 ( .DX(nn1854), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1000_), .F2(dummy_abc_1001_), .F3(dummy_abc_1002_) );
      defparam ii1854.CONFIG_DATA = 16'h5555;
      defparam ii1854.PLACE_LOCATION = "NONE";
      defparam ii1854.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1855 ( .DX(nn1855), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1003_), .F2(dummy_abc_1004_), .F3(dummy_abc_1005_) );
      defparam ii1855.CONFIG_DATA = 16'h5555;
      defparam ii1855.PLACE_LOCATION = "NONE";
      defparam ii1855.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1856 ( .DX(nn1856), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1006_), .F2(dummy_abc_1007_), .F3(dummy_abc_1008_) );
      defparam ii1856.CONFIG_DATA = 16'h5555;
      defparam ii1856.PLACE_LOCATION = "NONE";
      defparam ii1856.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1857 ( .DX(nn1857), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1009_), .F2(dummy_abc_1010_), .F3(dummy_abc_1011_) );
      defparam ii1857.CONFIG_DATA = 16'h5555;
      defparam ii1857.PLACE_LOCATION = "NONE";
      defparam ii1857.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1858 ( .DX(nn1858), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1012_), .F2(dummy_abc_1013_), .F3(dummy_abc_1014_) );
      defparam ii1858.CONFIG_DATA = 16'h5555;
      defparam ii1858.PLACE_LOCATION = "NONE";
      defparam ii1858.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1859 ( .DX(nn1859), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1015_), .F2(dummy_abc_1016_), .F3(dummy_abc_1017_) );
      defparam ii1859.CONFIG_DATA = 16'h5555;
      defparam ii1859.PLACE_LOCATION = "NONE";
      defparam ii1859.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1860 ( .DX(nn1860), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1018_), .F2(dummy_abc_1019_), .F3(dummy_abc_1020_) );
      defparam ii1860.CONFIG_DATA = 16'h5555;
      defparam ii1860.PLACE_LOCATION = "NONE";
      defparam ii1860.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1861 ( .DX(nn1861), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1021_), .F2(dummy_abc_1022_), .F3(dummy_abc_1023_) );
      defparam ii1861.CONFIG_DATA = 16'h5555;
      defparam ii1861.PLACE_LOCATION = "NONE";
      defparam ii1861.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1862 ( .DX(nn1862), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1024_), .F2(dummy_abc_1025_), .F3(dummy_abc_1026_) );
      defparam ii1862.CONFIG_DATA = 16'h5555;
      defparam ii1862.PLACE_LOCATION = "NONE";
      defparam ii1862.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1863 ( .DX(nn1863), .F0(dummy_abc_1027_), .F1(dummy_abc_1028_), .F2(dummy_abc_1029_), .F3(dummy_abc_1030_) );
      defparam ii1863.CONFIG_DATA = 16'hFFFF;
      defparam ii1863.PLACE_LOCATION = "NONE";
      defparam ii1863.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_265_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_622_ ), 
        .DX( {nn1863, nn1862, nn1861, nn1860, nn1859, nn1858, nn1857, nn1856, 
              nn1855, nn1854, nn1853, nn1852, nn1851, nn1850, nn1848, nn1846, 
              nn1844, nn1843} ), 
        .SUM( {\coefcal1_divide_inst2_u128_XORCI_17|SUM_net , dummy_623_, 
              dummy_624_, dummy_625_, dummy_626_, dummy_627_, dummy_628_, dummy_629_, 
              dummy_630_, dummy_631_, dummy_632_, dummy_633_, dummy_634_, dummy_635_, 
              dummy_636_, dummy_637_, dummy_638_, dummy_639_} )
      );
    CS_LUT4_PRIM ii1884 ( .DX(nn1884), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_603_), .F3(dummy_abc_1031_) );
      defparam ii1884.CONFIG_DATA = 16'hA6A6;
      defparam ii1884.PLACE_LOCATION = "NONE";
      defparam ii1884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1885 ( .DX(nn1885), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1032_), .F3(dummy_abc_1033_) );
      defparam ii1885.CONFIG_DATA = 16'h9999;
      defparam ii1885.PLACE_LOCATION = "NONE";
      defparam ii1885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1886 ( .DX(nn1886), .F0(\coefcal1_yDividend__reg[12]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_603_) );
      defparam ii1886.CONFIG_DATA = 16'hA569;
      defparam ii1886.PLACE_LOCATION = "NONE";
      defparam ii1886.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1887 ( .DX(nn1887), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn1845), .F2(dummy_abc_1034_), .F3(dummy_abc_1035_) );
      defparam ii1887.CONFIG_DATA = 16'h9999;
      defparam ii1887.PLACE_LOCATION = "NONE";
      defparam ii1887.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1888 ( .DX(nn1888), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1847), .F2(dummy_abc_1036_), .F3(dummy_abc_1037_) );
      defparam ii1888.CONFIG_DATA = 16'h9999;
      defparam ii1888.PLACE_LOCATION = "NONE";
      defparam ii1888.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1889 ( .DX(nn1889), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1849), .F2(dummy_abc_1038_), .F3(dummy_abc_1039_) );
      defparam ii1889.CONFIG_DATA = 16'h9999;
      defparam ii1889.PLACE_LOCATION = "NONE";
      defparam ii1889.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1890 ( .DX(nn1890), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1764), .F2(nn1842), .F3(dummy_abc_1040_) );
      defparam ii1890.CONFIG_DATA = 16'hD9D9;
      defparam ii1890.PLACE_LOCATION = "NONE";
      defparam ii1890.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1891 ( .DX(nn1891), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(dummy_abc_1041_), .F2(dummy_abc_1042_), .F3(dummy_abc_1043_) );
      defparam ii1891.CONFIG_DATA = 16'h5555;
      defparam ii1891.PLACE_LOCATION = "NONE";
      defparam ii1891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1892 ( .DX(nn1892), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_1044_), .F2(dummy_abc_1045_), .F3(dummy_abc_1046_) );
      defparam ii1892.CONFIG_DATA = 16'h5555;
      defparam ii1892.PLACE_LOCATION = "NONE";
      defparam ii1892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1893 ( .DX(nn1893), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1047_), .F2(dummy_abc_1048_), .F3(dummy_abc_1049_) );
      defparam ii1893.CONFIG_DATA = 16'h5555;
      defparam ii1893.PLACE_LOCATION = "NONE";
      defparam ii1893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1894 ( .DX(nn1894), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1050_), .F2(dummy_abc_1051_), .F3(dummy_abc_1052_) );
      defparam ii1894.CONFIG_DATA = 16'h5555;
      defparam ii1894.PLACE_LOCATION = "NONE";
      defparam ii1894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1895 ( .DX(nn1895), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1053_), .F2(dummy_abc_1054_), .F3(dummy_abc_1055_) );
      defparam ii1895.CONFIG_DATA = 16'h5555;
      defparam ii1895.PLACE_LOCATION = "NONE";
      defparam ii1895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1896 ( .DX(nn1896), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1056_), .F2(dummy_abc_1057_), .F3(dummy_abc_1058_) );
      defparam ii1896.CONFIG_DATA = 16'h5555;
      defparam ii1896.PLACE_LOCATION = "NONE";
      defparam ii1896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1897 ( .DX(nn1897), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1059_), .F2(dummy_abc_1060_), .F3(dummy_abc_1061_) );
      defparam ii1897.CONFIG_DATA = 16'h5555;
      defparam ii1897.PLACE_LOCATION = "NONE";
      defparam ii1897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1898 ( .DX(nn1898), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1062_), .F2(dummy_abc_1063_), .F3(dummy_abc_1064_) );
      defparam ii1898.CONFIG_DATA = 16'h5555;
      defparam ii1898.PLACE_LOCATION = "NONE";
      defparam ii1898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1899 ( .DX(nn1899), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1065_), .F2(dummy_abc_1066_), .F3(dummy_abc_1067_) );
      defparam ii1899.CONFIG_DATA = 16'h5555;
      defparam ii1899.PLACE_LOCATION = "NONE";
      defparam ii1899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1900 ( .DX(nn1900), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1068_), .F2(dummy_abc_1069_), .F3(dummy_abc_1070_) );
      defparam ii1900.CONFIG_DATA = 16'h5555;
      defparam ii1900.PLACE_LOCATION = "NONE";
      defparam ii1900.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1901 ( .DX(nn1901), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1071_), .F2(dummy_abc_1072_), .F3(dummy_abc_1073_) );
      defparam ii1901.CONFIG_DATA = 16'h5555;
      defparam ii1901.PLACE_LOCATION = "NONE";
      defparam ii1901.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_249_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn1849, nn1847, nn1845, nn1884, 
              \coefcal1_yDividend__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_179_ ), 
        .DX( {nn1901, nn1900, nn1899, nn1898, nn1897, nn1896, nn1895, nn1894, 
              nn1893, nn1892, nn1891, nn1890, nn1889, nn1888, nn1887, nn1886, 
              nn1885} ), 
        .SUM( {dummy_180_, \coefcal1_divide_inst2_u106_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_14|SUM_net , \coefcal1_divide_inst2_u106_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_12|SUM_net , \coefcal1_divide_inst2_u106_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_10|SUM_net , \coefcal1_divide_inst2_u106_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_8|SUM_net , \coefcal1_divide_inst2_u106_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_6|SUM_net , \coefcal1_divide_inst2_u106_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_4|SUM_net , \coefcal1_divide_inst2_u106_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_2|SUM_net , \coefcal1_divide_inst2_u106_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u106_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii1921 ( .DX(nn1921), .F0(nn1764), .F1(nn1842), .F2(dummy_622_), .F3(\coefcal1_divide_inst2_u106_XORCI_5|SUM_net ) );
      defparam ii1921.CONFIG_DATA = 16'h2A20;
      defparam ii1921.PLACE_LOCATION = "NONE";
      defparam ii1921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1922 ( .DX(nn1922), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1074_), .F3(dummy_abc_1075_) );
      defparam ii1922.CONFIG_DATA = 16'h9999;
      defparam ii1922.PLACE_LOCATION = "NONE";
      defparam ii1922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1923 ( .DX(nn1923), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_622_) );
      defparam ii1923.CONFIG_DATA = 16'hA569;
      defparam ii1923.PLACE_LOCATION = "NONE";
      defparam ii1923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1924 ( .DX(nn1924), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_622_), .F2(nn1884), .F3(\coefcal1_divide_inst2_u106_XORCI_1|SUM_net ) );
      defparam ii1924.CONFIG_DATA = 16'hA695;
      defparam ii1924.PLACE_LOCATION = "NONE";
      defparam ii1924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1925 ( .DX(nn1925), .F0(nn1845), .F1(dummy_622_), .F2(\coefcal1_divide_inst2_u106_XORCI_2|SUM_net ), .F3(dummy_abc_1076_) );
      defparam ii1925.CONFIG_DATA = 16'hB8B8;
      defparam ii1925.PLACE_LOCATION = "NONE";
      defparam ii1925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1926 ( .DX(nn1926), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1925), .F2(dummy_abc_1077_), .F3(dummy_abc_1078_) );
      defparam ii1926.CONFIG_DATA = 16'h9999;
      defparam ii1926.PLACE_LOCATION = "NONE";
      defparam ii1926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1927 ( .DX(nn1927), .F0(nn1847), .F1(dummy_622_), .F2(\coefcal1_divide_inst2_u106_XORCI_3|SUM_net ), .F3(dummy_abc_1079_) );
      defparam ii1927.CONFIG_DATA = 16'hB8B8;
      defparam ii1927.PLACE_LOCATION = "NONE";
      defparam ii1927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1928 ( .DX(nn1928), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1927), .F2(dummy_abc_1080_), .F3(dummy_abc_1081_) );
      defparam ii1928.CONFIG_DATA = 16'h9999;
      defparam ii1928.PLACE_LOCATION = "NONE";
      defparam ii1928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1929 ( .DX(nn1929), .F0(nn1849), .F1(dummy_622_), .F2(\coefcal1_divide_inst2_u106_XORCI_4|SUM_net ), .F3(dummy_abc_1082_) );
      defparam ii1929.CONFIG_DATA = 16'hB8B8;
      defparam ii1929.PLACE_LOCATION = "NONE";
      defparam ii1929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1930 ( .DX(nn1930), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1929), .F2(dummy_abc_1083_), .F3(dummy_abc_1084_) );
      defparam ii1930.CONFIG_DATA = 16'h9999;
      defparam ii1930.PLACE_LOCATION = "NONE";
      defparam ii1930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1931 ( .DX(nn1931), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1921), .F2(dummy_abc_1085_), .F3(dummy_abc_1086_) );
      defparam ii1931.CONFIG_DATA = 16'h9999;
      defparam ii1931.PLACE_LOCATION = "NONE";
      defparam ii1931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1932 ( .DX(nn1932), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_1087_), .F2(dummy_abc_1088_), .F3(dummy_abc_1089_) );
      defparam ii1932.CONFIG_DATA = 16'h5555;
      defparam ii1932.PLACE_LOCATION = "NONE";
      defparam ii1932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1933 ( .DX(nn1933), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1090_), .F2(dummy_abc_1091_), .F3(dummy_abc_1092_) );
      defparam ii1933.CONFIG_DATA = 16'h5555;
      defparam ii1933.PLACE_LOCATION = "NONE";
      defparam ii1933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1934 ( .DX(nn1934), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1093_), .F2(dummy_abc_1094_), .F3(dummy_abc_1095_) );
      defparam ii1934.CONFIG_DATA = 16'h5555;
      defparam ii1934.PLACE_LOCATION = "NONE";
      defparam ii1934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1935 ( .DX(nn1935), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1096_), .F2(dummy_abc_1097_), .F3(dummy_abc_1098_) );
      defparam ii1935.CONFIG_DATA = 16'h5555;
      defparam ii1935.PLACE_LOCATION = "NONE";
      defparam ii1935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1936 ( .DX(nn1936), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1099_), .F2(dummy_abc_1100_), .F3(dummy_abc_1101_) );
      defparam ii1936.CONFIG_DATA = 16'h5555;
      defparam ii1936.PLACE_LOCATION = "NONE";
      defparam ii1936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1937 ( .DX(nn1937), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1102_), .F2(dummy_abc_1103_), .F3(dummy_abc_1104_) );
      defparam ii1937.CONFIG_DATA = 16'h5555;
      defparam ii1937.PLACE_LOCATION = "NONE";
      defparam ii1937.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1938 ( .DX(nn1938), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1105_), .F2(dummy_abc_1106_), .F3(dummy_abc_1107_) );
      defparam ii1938.CONFIG_DATA = 16'h5555;
      defparam ii1938.PLACE_LOCATION = "NONE";
      defparam ii1938.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1939 ( .DX(nn1939), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1108_), .F2(dummy_abc_1109_), .F3(dummy_abc_1110_) );
      defparam ii1939.CONFIG_DATA = 16'h5555;
      defparam ii1939.PLACE_LOCATION = "NONE";
      defparam ii1939.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1940 ( .DX(nn1940), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1111_), .F2(dummy_abc_1112_), .F3(dummy_abc_1113_) );
      defparam ii1940.CONFIG_DATA = 16'h5555;
      defparam ii1940.PLACE_LOCATION = "NONE";
      defparam ii1940.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1941 ( .DX(nn1941), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1114_), .F2(dummy_abc_1115_), .F3(dummy_abc_1116_) );
      defparam ii1941.CONFIG_DATA = 16'h5555;
      defparam ii1941.PLACE_LOCATION = "NONE";
      defparam ii1941.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1942 ( .DX(nn1942), .F0(dummy_abc_1117_), .F1(dummy_abc_1118_), .F2(dummy_abc_1119_), .F3(dummy_abc_1120_) );
      defparam ii1942.CONFIG_DATA = 16'hFFFF;
      defparam ii1942.PLACE_LOCATION = "NONE";
      defparam ii1942.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_266_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_641_ ), 
        .DX( {nn1942, nn1941, nn1940, nn1939, nn1938, nn1937, nn1936, nn1935, 
              nn1934, nn1933, nn1932, nn1931, nn1930, nn1928, nn1926, nn1924, 
              nn1923, nn1922} ), 
        .SUM( {\coefcal1_divide_inst2_u130_XORCI_17|SUM_net , dummy_642_, 
              dummy_643_, dummy_644_, dummy_645_, dummy_646_, dummy_647_, dummy_648_, 
              dummy_649_, dummy_650_, dummy_651_, dummy_652_, dummy_653_, dummy_654_, 
              dummy_655_, dummy_656_, dummy_657_, dummy_658_} )
      );
    CS_LUT4_PRIM ii1963 ( .DX(nn1963), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1121_), .F3(dummy_abc_1122_) );
      defparam ii1963.CONFIG_DATA = 16'h9999;
      defparam ii1963.PLACE_LOCATION = "NONE";
      defparam ii1963.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1964 ( .DX(nn1964), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_641_) );
      defparam ii1964.CONFIG_DATA = 16'hA569;
      defparam ii1964.PLACE_LOCATION = "NONE";
      defparam ii1964.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1965 ( .DX(nn1965), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_622_), .F3(dummy_abc_1123_) );
      defparam ii1965.CONFIG_DATA = 16'hA6A6;
      defparam ii1965.PLACE_LOCATION = "NONE";
      defparam ii1965.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1966 ( .DX(nn1966), .F0(dummy_622_), .F1(nn1884), .F2(\coefcal1_divide_inst2_u106_XORCI_1|SUM_net ), .F3(dummy_abc_1124_) );
      defparam ii1966.CONFIG_DATA = 16'hD8D8;
      defparam ii1966.PLACE_LOCATION = "NONE";
      defparam ii1966.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1967 ( .DX(nn1967), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1125_), .F3(dummy_abc_1126_) );
      defparam ii1967.CONFIG_DATA = 16'h9999;
      defparam ii1967.PLACE_LOCATION = "NONE";
      defparam ii1967.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1968 ( .DX(nn1968), .F0(\coefcal1_yDividend__reg[11]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_622_) );
      defparam ii1968.CONFIG_DATA = 16'hA569;
      defparam ii1968.PLACE_LOCATION = "NONE";
      defparam ii1968.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1969 ( .DX(nn1969), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_622_), .F2(nn1884), .F3(\coefcal1_divide_inst2_u106_XORCI_1|SUM_net ) );
      defparam ii1969.CONFIG_DATA = 16'hA695;
      defparam ii1969.PLACE_LOCATION = "NONE";
      defparam ii1969.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1970 ( .DX(nn1970), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn1925), .F2(dummy_abc_1127_), .F3(dummy_abc_1128_) );
      defparam ii1970.CONFIG_DATA = 16'h9999;
      defparam ii1970.PLACE_LOCATION = "NONE";
      defparam ii1970.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1971 ( .DX(nn1971), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn1927), .F2(dummy_abc_1129_), .F3(dummy_abc_1130_) );
      defparam ii1971.CONFIG_DATA = 16'h9999;
      defparam ii1971.PLACE_LOCATION = "NONE";
      defparam ii1971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1972 ( .DX(nn1972), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn1929), .F2(dummy_abc_1131_), .F3(dummy_abc_1132_) );
      defparam ii1972.CONFIG_DATA = 16'h9999;
      defparam ii1972.PLACE_LOCATION = "NONE";
      defparam ii1972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1973 ( .DX(nn1973), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn1921), .F2(dummy_abc_1133_), .F3(dummy_abc_1134_) );
      defparam ii1973.CONFIG_DATA = 16'h9999;
      defparam ii1973.PLACE_LOCATION = "NONE";
      defparam ii1973.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1974 ( .DX(nn1974), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(dummy_abc_1135_), .F2(dummy_abc_1136_), .F3(dummy_abc_1137_) );
      defparam ii1974.CONFIG_DATA = 16'h5555;
      defparam ii1974.PLACE_LOCATION = "NONE";
      defparam ii1974.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1975 ( .DX(nn1975), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1138_), .F2(dummy_abc_1139_), .F3(dummy_abc_1140_) );
      defparam ii1975.CONFIG_DATA = 16'h5555;
      defparam ii1975.PLACE_LOCATION = "NONE";
      defparam ii1975.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1976 ( .DX(nn1976), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1141_), .F2(dummy_abc_1142_), .F3(dummy_abc_1143_) );
      defparam ii1976.CONFIG_DATA = 16'h5555;
      defparam ii1976.PLACE_LOCATION = "NONE";
      defparam ii1976.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1977 ( .DX(nn1977), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1144_), .F2(dummy_abc_1145_), .F3(dummy_abc_1146_) );
      defparam ii1977.CONFIG_DATA = 16'h5555;
      defparam ii1977.PLACE_LOCATION = "NONE";
      defparam ii1977.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1978 ( .DX(nn1978), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1147_), .F2(dummy_abc_1148_), .F3(dummy_abc_1149_) );
      defparam ii1978.CONFIG_DATA = 16'h5555;
      defparam ii1978.PLACE_LOCATION = "NONE";
      defparam ii1978.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1979 ( .DX(nn1979), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1150_), .F2(dummy_abc_1151_), .F3(dummy_abc_1152_) );
      defparam ii1979.CONFIG_DATA = 16'h5555;
      defparam ii1979.PLACE_LOCATION = "NONE";
      defparam ii1979.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1980 ( .DX(nn1980), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1153_), .F2(dummy_abc_1154_), .F3(dummy_abc_1155_) );
      defparam ii1980.CONFIG_DATA = 16'h5555;
      defparam ii1980.PLACE_LOCATION = "NONE";
      defparam ii1980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1981 ( .DX(nn1981), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1156_), .F2(dummy_abc_1157_), .F3(dummy_abc_1158_) );
      defparam ii1981.CONFIG_DATA = 16'h5555;
      defparam ii1981.PLACE_LOCATION = "NONE";
      defparam ii1981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1982 ( .DX(nn1982), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1159_), .F2(dummy_abc_1160_), .F3(dummy_abc_1161_) );
      defparam ii1982.CONFIG_DATA = 16'h5555;
      defparam ii1982.PLACE_LOCATION = "NONE";
      defparam ii1982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii1983 ( .DX(nn1983), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1162_), .F2(dummy_abc_1163_), .F3(dummy_abc_1164_) );
      defparam ii1983.CONFIG_DATA = 16'h5555;
      defparam ii1983.PLACE_LOCATION = "NONE";
      defparam ii1983.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_250_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn1921, nn1929, nn1927, nn1925, 
              nn1966, nn1965, \coefcal1_yDividend__reg[10]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_181_ ), 
        .DX( {nn1983, nn1982, nn1981, nn1980, nn1979, nn1978, nn1977, nn1976, 
              nn1975, nn1974, nn1973, nn1972, nn1971, nn1970, nn1969, nn1968, 
              nn1967} ), 
        .SUM( {dummy_182_, \coefcal1_divide_inst2_u107_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_14|SUM_net , \coefcal1_divide_inst2_u107_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_12|SUM_net , \coefcal1_divide_inst2_u107_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_10|SUM_net , \coefcal1_divide_inst2_u107_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_8|SUM_net , \coefcal1_divide_inst2_u107_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_6|SUM_net , \coefcal1_divide_inst2_u107_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_4|SUM_net , \coefcal1_divide_inst2_u107_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_2|SUM_net , \coefcal1_divide_inst2_u107_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u107_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2003 ( .DX(nn2003), .F0(dummy_641_), .F1(nn1965), .F2(\coefcal1_divide_inst2_u107_XORCI_1|SUM_net ), .F3(dummy_abc_1165_) );
      defparam ii2003.CONFIG_DATA = 16'hD8D8;
      defparam ii2003.PLACE_LOCATION = "NONE";
      defparam ii2003.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2004 ( .DX(nn2004), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2003), .F2(dummy_abc_1166_), .F3(dummy_abc_1167_) );
      defparam ii2004.CONFIG_DATA = 16'h9999;
      defparam ii2004.PLACE_LOCATION = "NONE";
      defparam ii2004.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2005 ( .DX(nn2005), .F0(nn1966), .F1(dummy_641_), .F2(\coefcal1_divide_inst2_u107_XORCI_2|SUM_net ), .F3(dummy_abc_1168_) );
      defparam ii2005.CONFIG_DATA = 16'hB8B8;
      defparam ii2005.PLACE_LOCATION = "NONE";
      defparam ii2005.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2006 ( .DX(nn2006), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2005), .F2(dummy_abc_1169_), .F3(dummy_abc_1170_) );
      defparam ii2006.CONFIG_DATA = 16'h9999;
      defparam ii2006.PLACE_LOCATION = "NONE";
      defparam ii2006.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2007 ( .DX(nn2007), .F0(nn1925), .F1(dummy_641_), .F2(\coefcal1_divide_inst2_u107_XORCI_3|SUM_net ), .F3(dummy_abc_1171_) );
      defparam ii2007.CONFIG_DATA = 16'hB8B8;
      defparam ii2007.PLACE_LOCATION = "NONE";
      defparam ii2007.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2008 ( .DX(nn2008), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2007), .F2(dummy_abc_1172_), .F3(dummy_abc_1173_) );
      defparam ii2008.CONFIG_DATA = 16'h9999;
      defparam ii2008.PLACE_LOCATION = "NONE";
      defparam ii2008.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2009 ( .DX(nn2009), .F0(nn1927), .F1(dummy_641_), .F2(\coefcal1_divide_inst2_u107_XORCI_4|SUM_net ), .F3(dummy_abc_1174_) );
      defparam ii2009.CONFIG_DATA = 16'hB8B8;
      defparam ii2009.PLACE_LOCATION = "NONE";
      defparam ii2009.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2010 ( .DX(nn2010), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2009), .F2(dummy_abc_1175_), .F3(dummy_abc_1176_) );
      defparam ii2010.CONFIG_DATA = 16'h9999;
      defparam ii2010.PLACE_LOCATION = "NONE";
      defparam ii2010.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2011 ( .DX(nn2011), .F0(nn1929), .F1(dummy_641_), .F2(\coefcal1_divide_inst2_u107_XORCI_5|SUM_net ), .F3(dummy_abc_1177_) );
      defparam ii2011.CONFIG_DATA = 16'hB8B8;
      defparam ii2011.PLACE_LOCATION = "NONE";
      defparam ii2011.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2012 ( .DX(nn2012), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2011), .F2(dummy_abc_1178_), .F3(dummy_abc_1179_) );
      defparam ii2012.CONFIG_DATA = 16'h9999;
      defparam ii2012.PLACE_LOCATION = "NONE";
      defparam ii2012.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2013 ( .DX(nn2013), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1921), .F2(dummy_641_), .F3(\coefcal1_divide_inst2_u107_XORCI_6|SUM_net ) );
      defparam ii2013.CONFIG_DATA = 16'h9A95;
      defparam ii2013.PLACE_LOCATION = "NONE";
      defparam ii2013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2014 ( .DX(nn2014), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1180_), .F2(dummy_abc_1181_), .F3(dummy_abc_1182_) );
      defparam ii2014.CONFIG_DATA = 16'h5555;
      defparam ii2014.PLACE_LOCATION = "NONE";
      defparam ii2014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2015 ( .DX(nn2015), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1183_), .F2(dummy_abc_1184_), .F3(dummy_abc_1185_) );
      defparam ii2015.CONFIG_DATA = 16'h5555;
      defparam ii2015.PLACE_LOCATION = "NONE";
      defparam ii2015.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2016 ( .DX(nn2016), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1186_), .F2(dummy_abc_1187_), .F3(dummy_abc_1188_) );
      defparam ii2016.CONFIG_DATA = 16'h5555;
      defparam ii2016.PLACE_LOCATION = "NONE";
      defparam ii2016.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2017 ( .DX(nn2017), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1189_), .F2(dummy_abc_1190_), .F3(dummy_abc_1191_) );
      defparam ii2017.CONFIG_DATA = 16'h5555;
      defparam ii2017.PLACE_LOCATION = "NONE";
      defparam ii2017.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2018 ( .DX(nn2018), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1192_), .F2(dummy_abc_1193_), .F3(dummy_abc_1194_) );
      defparam ii2018.CONFIG_DATA = 16'h5555;
      defparam ii2018.PLACE_LOCATION = "NONE";
      defparam ii2018.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2019 ( .DX(nn2019), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1195_), .F2(dummy_abc_1196_), .F3(dummy_abc_1197_) );
      defparam ii2019.CONFIG_DATA = 16'h5555;
      defparam ii2019.PLACE_LOCATION = "NONE";
      defparam ii2019.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2020 ( .DX(nn2020), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1198_), .F2(dummy_abc_1199_), .F3(dummy_abc_1200_) );
      defparam ii2020.CONFIG_DATA = 16'h5555;
      defparam ii2020.PLACE_LOCATION = "NONE";
      defparam ii2020.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2021 ( .DX(nn2021), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1201_), .F2(dummy_abc_1202_), .F3(dummy_abc_1203_) );
      defparam ii2021.CONFIG_DATA = 16'h5555;
      defparam ii2021.PLACE_LOCATION = "NONE";
      defparam ii2021.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2022 ( .DX(nn2022), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1204_), .F2(dummy_abc_1205_), .F3(dummy_abc_1206_) );
      defparam ii2022.CONFIG_DATA = 16'h5555;
      defparam ii2022.PLACE_LOCATION = "NONE";
      defparam ii2022.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2023 ( .DX(nn2023), .F0(dummy_abc_1207_), .F1(dummy_abc_1208_), .F2(dummy_abc_1209_), .F3(dummy_abc_1210_) );
      defparam ii2023.CONFIG_DATA = 16'hFFFF;
      defparam ii2023.PLACE_LOCATION = "NONE";
      defparam ii2023.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_267_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_660_ ), 
        .DX( {nn2023, nn2022, nn2021, nn2020, nn2019, nn2018, nn2017, nn2016, 
              nn2015, nn2014, nn2013, nn2012, nn2010, nn2008, nn2006, nn2004, 
              nn1964, nn1963} ), 
        .SUM( {\coefcal1_divide_inst2_u132_XORCI_17|SUM_net , dummy_661_, 
              dummy_662_, dummy_663_, dummy_664_, dummy_665_, dummy_666_, dummy_667_, 
              dummy_668_, dummy_669_, dummy_670_, dummy_671_, dummy_672_, dummy_673_, 
              dummy_674_, dummy_675_, dummy_676_, dummy_677_} )
      );
    CS_LUT4_PRIM ii2044 ( .DX(nn2044), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_641_), .F3(dummy_abc_1211_) );
      defparam ii2044.CONFIG_DATA = 16'hA6A6;
      defparam ii2044.PLACE_LOCATION = "NONE";
      defparam ii2044.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2045 ( .DX(nn2045), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1212_), .F3(dummy_abc_1213_) );
      defparam ii2045.CONFIG_DATA = 16'h9999;
      defparam ii2045.PLACE_LOCATION = "NONE";
      defparam ii2045.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2046 ( .DX(nn2046), .F0(\coefcal1_yDividend__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_641_) );
      defparam ii2046.CONFIG_DATA = 16'hA569;
      defparam ii2046.PLACE_LOCATION = "NONE";
      defparam ii2046.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2047 ( .DX(nn2047), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2003), .F2(dummy_abc_1214_), .F3(dummy_abc_1215_) );
      defparam ii2047.CONFIG_DATA = 16'h9999;
      defparam ii2047.PLACE_LOCATION = "NONE";
      defparam ii2047.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2048 ( .DX(nn2048), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2005), .F2(dummy_abc_1216_), .F3(dummy_abc_1217_) );
      defparam ii2048.CONFIG_DATA = 16'h9999;
      defparam ii2048.PLACE_LOCATION = "NONE";
      defparam ii2048.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2049 ( .DX(nn2049), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2007), .F2(dummy_abc_1218_), .F3(dummy_abc_1219_) );
      defparam ii2049.CONFIG_DATA = 16'h9999;
      defparam ii2049.PLACE_LOCATION = "NONE";
      defparam ii2049.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2050 ( .DX(nn2050), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2009), .F2(dummy_abc_1220_), .F3(dummy_abc_1221_) );
      defparam ii2050.CONFIG_DATA = 16'h9999;
      defparam ii2050.PLACE_LOCATION = "NONE";
      defparam ii2050.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2051 ( .DX(nn2051), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2011), .F2(dummy_abc_1222_), .F3(dummy_abc_1223_) );
      defparam ii2051.CONFIG_DATA = 16'h9999;
      defparam ii2051.PLACE_LOCATION = "NONE";
      defparam ii2051.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2052 ( .DX(nn2052), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn1921), .F2(dummy_641_), .F3(\coefcal1_divide_inst2_u107_XORCI_6|SUM_net ) );
      defparam ii2052.CONFIG_DATA = 16'h9A95;
      defparam ii2052.PLACE_LOCATION = "NONE";
      defparam ii2052.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2053 ( .DX(nn2053), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(dummy_abc_1224_), .F2(dummy_abc_1225_), .F3(dummy_abc_1226_) );
      defparam ii2053.CONFIG_DATA = 16'h5555;
      defparam ii2053.PLACE_LOCATION = "NONE";
      defparam ii2053.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2054 ( .DX(nn2054), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1227_), .F2(dummy_abc_1228_), .F3(dummy_abc_1229_) );
      defparam ii2054.CONFIG_DATA = 16'h5555;
      defparam ii2054.PLACE_LOCATION = "NONE";
      defparam ii2054.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2055 ( .DX(nn2055), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1230_), .F2(dummy_abc_1231_), .F3(dummy_abc_1232_) );
      defparam ii2055.CONFIG_DATA = 16'h5555;
      defparam ii2055.PLACE_LOCATION = "NONE";
      defparam ii2055.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2056 ( .DX(nn2056), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1233_), .F2(dummy_abc_1234_), .F3(dummy_abc_1235_) );
      defparam ii2056.CONFIG_DATA = 16'h5555;
      defparam ii2056.PLACE_LOCATION = "NONE";
      defparam ii2056.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2057 ( .DX(nn2057), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1236_), .F2(dummy_abc_1237_), .F3(dummy_abc_1238_) );
      defparam ii2057.CONFIG_DATA = 16'h5555;
      defparam ii2057.PLACE_LOCATION = "NONE";
      defparam ii2057.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2058 ( .DX(nn2058), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1239_), .F2(dummy_abc_1240_), .F3(dummy_abc_1241_) );
      defparam ii2058.CONFIG_DATA = 16'h5555;
      defparam ii2058.PLACE_LOCATION = "NONE";
      defparam ii2058.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2059 ( .DX(nn2059), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1242_), .F2(dummy_abc_1243_), .F3(dummy_abc_1244_) );
      defparam ii2059.CONFIG_DATA = 16'h5555;
      defparam ii2059.PLACE_LOCATION = "NONE";
      defparam ii2059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2060 ( .DX(nn2060), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1245_), .F2(dummy_abc_1246_), .F3(dummy_abc_1247_) );
      defparam ii2060.CONFIG_DATA = 16'h5555;
      defparam ii2060.PLACE_LOCATION = "NONE";
      defparam ii2060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2061 ( .DX(nn2061), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1248_), .F2(dummy_abc_1249_), .F3(dummy_abc_1250_) );
      defparam ii2061.CONFIG_DATA = 16'h5555;
      defparam ii2061.PLACE_LOCATION = "NONE";
      defparam ii2061.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_251_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, 1'b0, nn2011, nn2009, nn2007, nn2005, nn2003, nn2044, 
              \coefcal1_yDividend__reg[9]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_183_ ), 
        .DX( {nn2061, nn2060, nn2059, nn2058, nn2057, nn2056, nn2055, nn2054, 
              nn2053, nn2052, nn2051, nn2050, nn2049, nn2048, nn2047, nn2046, 
              nn2045} ), 
        .SUM( {dummy_184_, \coefcal1_divide_inst2_u108_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_14|SUM_net , \coefcal1_divide_inst2_u108_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_12|SUM_net , \coefcal1_divide_inst2_u108_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_10|SUM_net , \coefcal1_divide_inst2_u108_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_8|SUM_net , \coefcal1_divide_inst2_u108_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_6|SUM_net , \coefcal1_divide_inst2_u108_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_4|SUM_net , \coefcal1_divide_inst2_u108_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_2|SUM_net , \coefcal1_divide_inst2_u108_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2081 ( .DX(nn2081), .F0(nn1921), .F1(dummy_641_), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ) );
      defparam ii2081.CONFIG_DATA = 16'h8F80;
      defparam ii2081.PLACE_LOCATION = "NONE";
      defparam ii2081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2082 ( .DX(nn2082), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1251_), .F3(dummy_abc_1252_) );
      defparam ii2082.CONFIG_DATA = 16'h9999;
      defparam ii2082.PLACE_LOCATION = "NONE";
      defparam ii2082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2083 ( .DX(nn2083), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_660_) );
      defparam ii2083.CONFIG_DATA = 16'hA569;
      defparam ii2083.PLACE_LOCATION = "NONE";
      defparam ii2083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2084 ( .DX(nn2084), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_660_), .F2(nn2044), .F3(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ) );
      defparam ii2084.CONFIG_DATA = 16'hA695;
      defparam ii2084.PLACE_LOCATION = "NONE";
      defparam ii2084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2085 ( .DX(nn2085), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2003), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ) );
      defparam ii2085.CONFIG_DATA = 16'h9A95;
      defparam ii2085.PLACE_LOCATION = "NONE";
      defparam ii2085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2086 ( .DX(nn2086), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2005), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ) );
      defparam ii2086.CONFIG_DATA = 16'h9A95;
      defparam ii2086.PLACE_LOCATION = "NONE";
      defparam ii2086.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2087 ( .DX(nn2087), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2007), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ) );
      defparam ii2087.CONFIG_DATA = 16'h9A95;
      defparam ii2087.PLACE_LOCATION = "NONE";
      defparam ii2087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2088 ( .DX(nn2088), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2009), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ) );
      defparam ii2088.CONFIG_DATA = 16'h9A95;
      defparam ii2088.PLACE_LOCATION = "NONE";
      defparam ii2088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2089 ( .DX(nn2089), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2011), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ) );
      defparam ii2089.CONFIG_DATA = 16'h9A95;
      defparam ii2089.PLACE_LOCATION = "NONE";
      defparam ii2089.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2090 ( .DX(nn2090), .F0(nn1921), .F1(dummy_641_), .F2(dummy_abc_1253_), .F3(dummy_abc_1254_) );
      defparam ii2090.CONFIG_DATA = 16'h8888;
      defparam ii2090.PLACE_LOCATION = "NONE";
      defparam ii2090.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2091 ( .DX(nn2091), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2090), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ) );
      defparam ii2091.CONFIG_DATA = 16'h9095;
      defparam ii2091.PLACE_LOCATION = "NONE";
      defparam ii2091.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2092 ( .DX(nn2092), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1255_), .F2(dummy_abc_1256_), .F3(dummy_abc_1257_) );
      defparam ii2092.CONFIG_DATA = 16'h5555;
      defparam ii2092.PLACE_LOCATION = "NONE";
      defparam ii2092.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2093 ( .DX(nn2093), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1258_), .F2(dummy_abc_1259_), .F3(dummy_abc_1260_) );
      defparam ii2093.CONFIG_DATA = 16'h5555;
      defparam ii2093.PLACE_LOCATION = "NONE";
      defparam ii2093.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2094 ( .DX(nn2094), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1261_), .F2(dummy_abc_1262_), .F3(dummy_abc_1263_) );
      defparam ii2094.CONFIG_DATA = 16'h5555;
      defparam ii2094.PLACE_LOCATION = "NONE";
      defparam ii2094.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2095 ( .DX(nn2095), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1264_), .F2(dummy_abc_1265_), .F3(dummy_abc_1266_) );
      defparam ii2095.CONFIG_DATA = 16'h5555;
      defparam ii2095.PLACE_LOCATION = "NONE";
      defparam ii2095.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2096 ( .DX(nn2096), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1267_), .F2(dummy_abc_1268_), .F3(dummy_abc_1269_) );
      defparam ii2096.CONFIG_DATA = 16'h5555;
      defparam ii2096.PLACE_LOCATION = "NONE";
      defparam ii2096.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2097 ( .DX(nn2097), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1270_), .F2(dummy_abc_1271_), .F3(dummy_abc_1272_) );
      defparam ii2097.CONFIG_DATA = 16'h5555;
      defparam ii2097.PLACE_LOCATION = "NONE";
      defparam ii2097.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2098 ( .DX(nn2098), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1273_), .F2(dummy_abc_1274_), .F3(dummy_abc_1275_) );
      defparam ii2098.CONFIG_DATA = 16'h5555;
      defparam ii2098.PLACE_LOCATION = "NONE";
      defparam ii2098.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2099 ( .DX(nn2099), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1276_), .F2(dummy_abc_1277_), .F3(dummy_abc_1278_) );
      defparam ii2099.CONFIG_DATA = 16'h5555;
      defparam ii2099.PLACE_LOCATION = "NONE";
      defparam ii2099.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2100 ( .DX(nn2100), .F0(dummy_abc_1279_), .F1(dummy_abc_1280_), .F2(dummy_abc_1281_), .F3(dummy_abc_1282_) );
      defparam ii2100.CONFIG_DATA = 16'hFFFF;
      defparam ii2100.PLACE_LOCATION = "NONE";
      defparam ii2100.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_268_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_679_ ), 
        .DX( {nn2100, nn2099, nn2098, nn2097, nn2096, nn2095, nn2094, nn2093, 
              nn2092, nn2091, nn2089, nn2088, nn2087, nn2086, nn2085, nn2084, 
              nn2083, nn2082} ), 
        .SUM( {\coefcal1_divide_inst2_u134_XORCI_17|SUM_net , dummy_680_, 
              dummy_681_, dummy_682_, dummy_683_, dummy_684_, dummy_685_, dummy_686_, 
              dummy_687_, dummy_688_, dummy_689_, dummy_690_, dummy_691_, dummy_692_, 
              dummy_693_, dummy_694_, dummy_695_, dummy_696_} )
      );
    CS_LUT4_PRIM ii2121 ( .DX(nn2121), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_660_), .F3(dummy_abc_1283_) );
      defparam ii2121.CONFIG_DATA = 16'hA6A6;
      defparam ii2121.PLACE_LOCATION = "NONE";
      defparam ii2121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2122 ( .DX(nn2122), .F0(dummy_660_), .F1(nn2044), .F2(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ), .F3(dummy_abc_1284_) );
      defparam ii2122.CONFIG_DATA = 16'hD8D8;
      defparam ii2122.PLACE_LOCATION = "NONE";
      defparam ii2122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2123 ( .DX(nn2123), .F0(nn2003), .F1(dummy_660_), .F2(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ), .F3(dummy_abc_1285_) );
      defparam ii2123.CONFIG_DATA = 16'hB8B8;
      defparam ii2123.PLACE_LOCATION = "NONE";
      defparam ii2123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2124 ( .DX(nn2124), .F0(nn2005), .F1(dummy_660_), .F2(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ), .F3(dummy_abc_1286_) );
      defparam ii2124.CONFIG_DATA = 16'hB8B8;
      defparam ii2124.PLACE_LOCATION = "NONE";
      defparam ii2124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2125 ( .DX(nn2125), .F0(nn2007), .F1(dummy_660_), .F2(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ), .F3(dummy_abc_1287_) );
      defparam ii2125.CONFIG_DATA = 16'hB8B8;
      defparam ii2125.PLACE_LOCATION = "NONE";
      defparam ii2125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2126 ( .DX(nn2126), .F0(nn2009), .F1(dummy_660_), .F2(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ), .F3(dummy_abc_1288_) );
      defparam ii2126.CONFIG_DATA = 16'hB8B8;
      defparam ii2126.PLACE_LOCATION = "NONE";
      defparam ii2126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2127 ( .DX(nn2127), .F0(nn2011), .F1(dummy_660_), .F2(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ), .F3(dummy_abc_1289_) );
      defparam ii2127.CONFIG_DATA = 16'hB8B8;
      defparam ii2127.PLACE_LOCATION = "NONE";
      defparam ii2127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2128 ( .DX(nn2128), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1290_), .F3(dummy_abc_1291_) );
      defparam ii2128.CONFIG_DATA = 16'h9999;
      defparam ii2128.PLACE_LOCATION = "NONE";
      defparam ii2128.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2129 ( .DX(nn2129), .F0(\coefcal1_yDividend__reg[9]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_660_) );
      defparam ii2129.CONFIG_DATA = 16'hA569;
      defparam ii2129.PLACE_LOCATION = "NONE";
      defparam ii2129.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2130 ( .DX(nn2130), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_660_), .F2(nn2044), .F3(\coefcal1_divide_inst2_u108_XORCI_1|SUM_net ) );
      defparam ii2130.CONFIG_DATA = 16'hA695;
      defparam ii2130.PLACE_LOCATION = "NONE";
      defparam ii2130.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2131 ( .DX(nn2131), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2003), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_2|SUM_net ) );
      defparam ii2131.CONFIG_DATA = 16'h9A95;
      defparam ii2131.PLACE_LOCATION = "NONE";
      defparam ii2131.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2132 ( .DX(nn2132), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2005), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_3|SUM_net ) );
      defparam ii2132.CONFIG_DATA = 16'h9A95;
      defparam ii2132.PLACE_LOCATION = "NONE";
      defparam ii2132.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2133 ( .DX(nn2133), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2007), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_4|SUM_net ) );
      defparam ii2133.CONFIG_DATA = 16'h9A95;
      defparam ii2133.PLACE_LOCATION = "NONE";
      defparam ii2133.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2134 ( .DX(nn2134), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2009), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_5|SUM_net ) );
      defparam ii2134.CONFIG_DATA = 16'h9A95;
      defparam ii2134.PLACE_LOCATION = "NONE";
      defparam ii2134.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2135 ( .DX(nn2135), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2011), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_6|SUM_net ) );
      defparam ii2135.CONFIG_DATA = 16'h9A95;
      defparam ii2135.PLACE_LOCATION = "NONE";
      defparam ii2135.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2136 ( .DX(nn2136), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2090), .F2(dummy_660_), .F3(\coefcal1_divide_inst2_u108_XORCI_7|SUM_net ) );
      defparam ii2136.CONFIG_DATA = 16'h9095;
      defparam ii2136.PLACE_LOCATION = "NONE";
      defparam ii2136.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2137 ( .DX(nn2137), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(dummy_abc_1292_), .F2(dummy_abc_1293_), .F3(dummy_abc_1294_) );
      defparam ii2137.CONFIG_DATA = 16'h5555;
      defparam ii2137.PLACE_LOCATION = "NONE";
      defparam ii2137.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2138 ( .DX(nn2138), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1295_), .F2(dummy_abc_1296_), .F3(dummy_abc_1297_) );
      defparam ii2138.CONFIG_DATA = 16'h5555;
      defparam ii2138.PLACE_LOCATION = "NONE";
      defparam ii2138.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2139 ( .DX(nn2139), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1298_), .F2(dummy_abc_1299_), .F3(dummy_abc_1300_) );
      defparam ii2139.CONFIG_DATA = 16'h5555;
      defparam ii2139.PLACE_LOCATION = "NONE";
      defparam ii2139.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2140 ( .DX(nn2140), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1301_), .F2(dummy_abc_1302_), .F3(dummy_abc_1303_) );
      defparam ii2140.CONFIG_DATA = 16'h5555;
      defparam ii2140.PLACE_LOCATION = "NONE";
      defparam ii2140.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2141 ( .DX(nn2141), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1304_), .F2(dummy_abc_1305_), .F3(dummy_abc_1306_) );
      defparam ii2141.CONFIG_DATA = 16'h5555;
      defparam ii2141.PLACE_LOCATION = "NONE";
      defparam ii2141.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2142 ( .DX(nn2142), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1307_), .F2(dummy_abc_1308_), .F3(dummy_abc_1309_) );
      defparam ii2142.CONFIG_DATA = 16'h5555;
      defparam ii2142.PLACE_LOCATION = "NONE";
      defparam ii2142.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2143 ( .DX(nn2143), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1310_), .F2(dummy_abc_1311_), .F3(dummy_abc_1312_) );
      defparam ii2143.CONFIG_DATA = 16'h5555;
      defparam ii2143.PLACE_LOCATION = "NONE";
      defparam ii2143.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2144 ( .DX(nn2144), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1313_), .F2(dummy_abc_1314_), .F3(dummy_abc_1315_) );
      defparam ii2144.CONFIG_DATA = 16'h5555;
      defparam ii2144.PLACE_LOCATION = "NONE";
      defparam ii2144.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_252_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn2081, 
              nn2127, nn2126, nn2125, nn2124, nn2123, nn2122, nn2121, 
              \coefcal1_yDividend__reg[8]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_185_ ), 
        .DX( {nn2144, nn2143, nn2142, nn2141, nn2140, nn2139, nn2138, nn2137, 
              nn2136, nn2135, nn2134, nn2133, nn2132, nn2131, nn2130, nn2129, 
              nn2128} ), 
        .SUM( {dummy_186_, \coefcal1_divide_inst2_u109_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_14|SUM_net , \coefcal1_divide_inst2_u109_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_12|SUM_net , \coefcal1_divide_inst2_u109_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_10|SUM_net , \coefcal1_divide_inst2_u109_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_8|SUM_net , \coefcal1_divide_inst2_u109_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_6|SUM_net , \coefcal1_divide_inst2_u109_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_4|SUM_net , \coefcal1_divide_inst2_u109_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_2|SUM_net , \coefcal1_divide_inst2_u109_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u109_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2164 ( .DX(nn2164), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1316_), .F3(dummy_abc_1317_) );
      defparam ii2164.CONFIG_DATA = 16'h9999;
      defparam ii2164.PLACE_LOCATION = "NONE";
      defparam ii2164.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2165 ( .DX(nn2165), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_679_) );
      defparam ii2165.CONFIG_DATA = 16'hA569;
      defparam ii2165.PLACE_LOCATION = "NONE";
      defparam ii2165.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2166 ( .DX(nn2166), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_679_), .F2(nn2121), .F3(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ) );
      defparam ii2166.CONFIG_DATA = 16'hA695;
      defparam ii2166.PLACE_LOCATION = "NONE";
      defparam ii2166.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2167 ( .DX(nn2167), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2122), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ) );
      defparam ii2167.CONFIG_DATA = 16'h9A95;
      defparam ii2167.PLACE_LOCATION = "NONE";
      defparam ii2167.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2168 ( .DX(nn2168), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2123), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ) );
      defparam ii2168.CONFIG_DATA = 16'h9A95;
      defparam ii2168.PLACE_LOCATION = "NONE";
      defparam ii2168.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2169 ( .DX(nn2169), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2124), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ) );
      defparam ii2169.CONFIG_DATA = 16'h9A95;
      defparam ii2169.PLACE_LOCATION = "NONE";
      defparam ii2169.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2170 ( .DX(nn2170), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2125), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ) );
      defparam ii2170.CONFIG_DATA = 16'h9A95;
      defparam ii2170.PLACE_LOCATION = "NONE";
      defparam ii2170.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2171 ( .DX(nn2171), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2126), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ) );
      defparam ii2171.CONFIG_DATA = 16'h9A95;
      defparam ii2171.PLACE_LOCATION = "NONE";
      defparam ii2171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2172 ( .DX(nn2172), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2127), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ) );
      defparam ii2172.CONFIG_DATA = 16'h9A95;
      defparam ii2172.PLACE_LOCATION = "NONE";
      defparam ii2172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2173 ( .DX(nn2173), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2081), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ) );
      defparam ii2173.CONFIG_DATA = 16'h9995;
      defparam ii2173.PLACE_LOCATION = "NONE";
      defparam ii2173.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2174 ( .DX(nn2174), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1318_), .F2(dummy_abc_1319_), .F3(dummy_abc_1320_) );
      defparam ii2174.CONFIG_DATA = 16'h5555;
      defparam ii2174.PLACE_LOCATION = "NONE";
      defparam ii2174.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2175 ( .DX(nn2175), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1321_), .F2(dummy_abc_1322_), .F3(dummy_abc_1323_) );
      defparam ii2175.CONFIG_DATA = 16'h5555;
      defparam ii2175.PLACE_LOCATION = "NONE";
      defparam ii2175.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2176 ( .DX(nn2176), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1324_), .F2(dummy_abc_1325_), .F3(dummy_abc_1326_) );
      defparam ii2176.CONFIG_DATA = 16'h5555;
      defparam ii2176.PLACE_LOCATION = "NONE";
      defparam ii2176.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2177 ( .DX(nn2177), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1327_), .F2(dummy_abc_1328_), .F3(dummy_abc_1329_) );
      defparam ii2177.CONFIG_DATA = 16'h5555;
      defparam ii2177.PLACE_LOCATION = "NONE";
      defparam ii2177.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2178 ( .DX(nn2178), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1330_), .F2(dummy_abc_1331_), .F3(dummy_abc_1332_) );
      defparam ii2178.CONFIG_DATA = 16'h5555;
      defparam ii2178.PLACE_LOCATION = "NONE";
      defparam ii2178.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2179 ( .DX(nn2179), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1333_), .F2(dummy_abc_1334_), .F3(dummy_abc_1335_) );
      defparam ii2179.CONFIG_DATA = 16'h5555;
      defparam ii2179.PLACE_LOCATION = "NONE";
      defparam ii2179.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2180 ( .DX(nn2180), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1336_), .F2(dummy_abc_1337_), .F3(dummy_abc_1338_) );
      defparam ii2180.CONFIG_DATA = 16'h5555;
      defparam ii2180.PLACE_LOCATION = "NONE";
      defparam ii2180.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2181 ( .DX(nn2181), .F0(dummy_abc_1339_), .F1(dummy_abc_1340_), .F2(dummy_abc_1341_), .F3(dummy_abc_1342_) );
      defparam ii2181.CONFIG_DATA = 16'hFFFF;
      defparam ii2181.PLACE_LOCATION = "NONE";
      defparam ii2181.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_269_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_698_ ), 
        .DX( {nn2181, nn2180, nn2179, nn2178, nn2177, nn2176, nn2175, nn2174, 
              nn2173, nn2172, nn2171, nn2170, nn2169, nn2168, nn2167, nn2166, 
              nn2165, nn2164} ), 
        .SUM( {\coefcal1_divide_inst2_u136_XORCI_17|SUM_net , dummy_699_, 
              dummy_700_, dummy_701_, dummy_702_, dummy_703_, dummy_704_, dummy_705_, 
              dummy_706_, dummy_707_, dummy_708_, dummy_709_, dummy_710_, dummy_711_, 
              dummy_712_, dummy_713_, dummy_714_, dummy_715_} )
      );
    CS_LUT4_PRIM ii2202 ( .DX(nn2202), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_679_), .F3(dummy_abc_1343_) );
      defparam ii2202.CONFIG_DATA = 16'hA6A6;
      defparam ii2202.PLACE_LOCATION = "NONE";
      defparam ii2202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2203 ( .DX(nn2203), .F0(dummy_679_), .F1(nn2121), .F2(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ), .F3(dummy_abc_1344_) );
      defparam ii2203.CONFIG_DATA = 16'hD8D8;
      defparam ii2203.PLACE_LOCATION = "NONE";
      defparam ii2203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2204 ( .DX(nn2204), .F0(nn2122), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ), .F3(dummy_abc_1345_) );
      defparam ii2204.CONFIG_DATA = 16'hB8B8;
      defparam ii2204.PLACE_LOCATION = "NONE";
      defparam ii2204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2205 ( .DX(nn2205), .F0(nn2123), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ), .F3(dummy_abc_1346_) );
      defparam ii2205.CONFIG_DATA = 16'hB8B8;
      defparam ii2205.PLACE_LOCATION = "NONE";
      defparam ii2205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2206 ( .DX(nn2206), .F0(nn2124), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ), .F3(dummy_abc_1347_) );
      defparam ii2206.CONFIG_DATA = 16'hB8B8;
      defparam ii2206.PLACE_LOCATION = "NONE";
      defparam ii2206.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2207 ( .DX(nn2207), .F0(nn2125), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ), .F3(dummy_abc_1348_) );
      defparam ii2207.CONFIG_DATA = 16'hB8B8;
      defparam ii2207.PLACE_LOCATION = "NONE";
      defparam ii2207.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2208 ( .DX(nn2208), .F0(nn2126), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ), .F3(dummy_abc_1349_) );
      defparam ii2208.CONFIG_DATA = 16'hB8B8;
      defparam ii2208.PLACE_LOCATION = "NONE";
      defparam ii2208.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2209 ( .DX(nn2209), .F0(nn2127), .F1(dummy_679_), .F2(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ), .F3(dummy_abc_1350_) );
      defparam ii2209.CONFIG_DATA = 16'hB8B8;
      defparam ii2209.PLACE_LOCATION = "NONE";
      defparam ii2209.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2210 ( .DX(nn2210), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1351_), .F3(dummy_abc_1352_) );
      defparam ii2210.CONFIG_DATA = 16'h9999;
      defparam ii2210.PLACE_LOCATION = "NONE";
      defparam ii2210.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2211 ( .DX(nn2211), .F0(\coefcal1_yDividend__reg[8]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_679_) );
      defparam ii2211.CONFIG_DATA = 16'hA569;
      defparam ii2211.PLACE_LOCATION = "NONE";
      defparam ii2211.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2212 ( .DX(nn2212), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_679_), .F2(nn2121), .F3(\coefcal1_divide_inst2_u109_XORCI_1|SUM_net ) );
      defparam ii2212.CONFIG_DATA = 16'hA695;
      defparam ii2212.PLACE_LOCATION = "NONE";
      defparam ii2212.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2213 ( .DX(nn2213), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2122), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_2|SUM_net ) );
      defparam ii2213.CONFIG_DATA = 16'h9A95;
      defparam ii2213.PLACE_LOCATION = "NONE";
      defparam ii2213.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2214 ( .DX(nn2214), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2123), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_3|SUM_net ) );
      defparam ii2214.CONFIG_DATA = 16'h9A95;
      defparam ii2214.PLACE_LOCATION = "NONE";
      defparam ii2214.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2215 ( .DX(nn2215), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2124), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_4|SUM_net ) );
      defparam ii2215.CONFIG_DATA = 16'h9A95;
      defparam ii2215.PLACE_LOCATION = "NONE";
      defparam ii2215.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2216 ( .DX(nn2216), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2125), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_5|SUM_net ) );
      defparam ii2216.CONFIG_DATA = 16'h9A95;
      defparam ii2216.PLACE_LOCATION = "NONE";
      defparam ii2216.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2217 ( .DX(nn2217), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2126), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_6|SUM_net ) );
      defparam ii2217.CONFIG_DATA = 16'h9A95;
      defparam ii2217.PLACE_LOCATION = "NONE";
      defparam ii2217.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2218 ( .DX(nn2218), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2127), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_7|SUM_net ) );
      defparam ii2218.CONFIG_DATA = 16'h9A95;
      defparam ii2218.PLACE_LOCATION = "NONE";
      defparam ii2218.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2219 ( .DX(nn2219), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2081), .F2(dummy_679_), .F3(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ) );
      defparam ii2219.CONFIG_DATA = 16'h9995;
      defparam ii2219.PLACE_LOCATION = "NONE";
      defparam ii2219.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2220 ( .DX(nn2220), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(dummy_abc_1353_), .F2(dummy_abc_1354_), .F3(dummy_abc_1355_) );
      defparam ii2220.CONFIG_DATA = 16'h5555;
      defparam ii2220.PLACE_LOCATION = "NONE";
      defparam ii2220.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2221 ( .DX(nn2221), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1356_), .F2(dummy_abc_1357_), .F3(dummy_abc_1358_) );
      defparam ii2221.CONFIG_DATA = 16'h5555;
      defparam ii2221.PLACE_LOCATION = "NONE";
      defparam ii2221.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2222 ( .DX(nn2222), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1359_), .F2(dummy_abc_1360_), .F3(dummy_abc_1361_) );
      defparam ii2222.CONFIG_DATA = 16'h5555;
      defparam ii2222.PLACE_LOCATION = "NONE";
      defparam ii2222.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2223 ( .DX(nn2223), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1362_), .F2(dummy_abc_1363_), .F3(dummy_abc_1364_) );
      defparam ii2223.CONFIG_DATA = 16'h5555;
      defparam ii2223.PLACE_LOCATION = "NONE";
      defparam ii2223.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2224 ( .DX(nn2224), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1365_), .F2(dummy_abc_1366_), .F3(dummy_abc_1367_) );
      defparam ii2224.CONFIG_DATA = 16'h5555;
      defparam ii2224.PLACE_LOCATION = "NONE";
      defparam ii2224.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2225 ( .DX(nn2225), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1368_), .F2(dummy_abc_1369_), .F3(dummy_abc_1370_) );
      defparam ii2225.CONFIG_DATA = 16'h5555;
      defparam ii2225.PLACE_LOCATION = "NONE";
      defparam ii2225.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2226 ( .DX(nn2226), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1371_), .F2(dummy_abc_1372_), .F3(dummy_abc_1373_) );
      defparam ii2226.CONFIG_DATA = 16'h5555;
      defparam ii2226.PLACE_LOCATION = "NONE";
      defparam ii2226.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_253_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn2209, 
              nn2208, nn2207, nn2206, nn2205, nn2204, nn2203, nn2202, 
              \coefcal1_yDividend__reg[7]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_187_ ), 
        .DX( {nn2226, nn2225, nn2224, nn2223, nn2222, nn2221, nn2220, nn2219, 
              nn2218, nn2217, nn2216, nn2215, nn2214, nn2213, nn2212, nn2211, 
              nn2210} ), 
        .SUM( {dummy_188_, \coefcal1_divide_inst2_u110_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_14|SUM_net , \coefcal1_divide_inst2_u110_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_12|SUM_net , \coefcal1_divide_inst2_u110_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_10|SUM_net , \coefcal1_divide_inst2_u110_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_8|SUM_net , \coefcal1_divide_inst2_u110_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_6|SUM_net , \coefcal1_divide_inst2_u110_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_4|SUM_net , \coefcal1_divide_inst2_u110_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_2|SUM_net , \coefcal1_divide_inst2_u110_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2246 ( .DX(nn2246), .F0(dummy_679_), .F1(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ), .F2(dummy_698_), .F3(\coefcal1_divide_inst2_u110_XORCI_9|SUM_net ) );
      defparam ii2246.CONFIG_DATA = 16'hEFE0;
      defparam ii2246.PLACE_LOCATION = "NONE";
      defparam ii2246.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2247 ( .DX(nn2247), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1374_), .F3(dummy_abc_1375_) );
      defparam ii2247.CONFIG_DATA = 16'h9999;
      defparam ii2247.PLACE_LOCATION = "NONE";
      defparam ii2247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2248 ( .DX(nn2248), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_698_) );
      defparam ii2248.CONFIG_DATA = 16'hA569;
      defparam ii2248.PLACE_LOCATION = "NONE";
      defparam ii2248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2249 ( .DX(nn2249), .F0(dummy_698_), .F1(nn2202), .F2(\coefcal1_divide_inst2_u110_XORCI_1|SUM_net ), .F3(dummy_abc_1376_) );
      defparam ii2249.CONFIG_DATA = 16'hD8D8;
      defparam ii2249.PLACE_LOCATION = "NONE";
      defparam ii2249.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2250 ( .DX(nn2250), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2249), .F2(dummy_abc_1377_), .F3(dummy_abc_1378_) );
      defparam ii2250.CONFIG_DATA = 16'h9999;
      defparam ii2250.PLACE_LOCATION = "NONE";
      defparam ii2250.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2251 ( .DX(nn2251), .F0(nn2203), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_2|SUM_net ), .F3(dummy_abc_1379_) );
      defparam ii2251.CONFIG_DATA = 16'hB8B8;
      defparam ii2251.PLACE_LOCATION = "NONE";
      defparam ii2251.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2252 ( .DX(nn2252), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2251), .F2(dummy_abc_1380_), .F3(dummy_abc_1381_) );
      defparam ii2252.CONFIG_DATA = 16'h9999;
      defparam ii2252.PLACE_LOCATION = "NONE";
      defparam ii2252.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2253 ( .DX(nn2253), .F0(nn2204), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_3|SUM_net ), .F3(dummy_abc_1382_) );
      defparam ii2253.CONFIG_DATA = 16'hB8B8;
      defparam ii2253.PLACE_LOCATION = "NONE";
      defparam ii2253.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2254 ( .DX(nn2254), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2253), .F2(dummy_abc_1383_), .F3(dummy_abc_1384_) );
      defparam ii2254.CONFIG_DATA = 16'h9999;
      defparam ii2254.PLACE_LOCATION = "NONE";
      defparam ii2254.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2255 ( .DX(nn2255), .F0(nn2205), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_4|SUM_net ), .F3(dummy_abc_1385_) );
      defparam ii2255.CONFIG_DATA = 16'hB8B8;
      defparam ii2255.PLACE_LOCATION = "NONE";
      defparam ii2255.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2256 ( .DX(nn2256), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2255), .F2(dummy_abc_1386_), .F3(dummy_abc_1387_) );
      defparam ii2256.CONFIG_DATA = 16'h9999;
      defparam ii2256.PLACE_LOCATION = "NONE";
      defparam ii2256.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2257 ( .DX(nn2257), .F0(nn2206), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_5|SUM_net ), .F3(dummy_abc_1388_) );
      defparam ii2257.CONFIG_DATA = 16'hB8B8;
      defparam ii2257.PLACE_LOCATION = "NONE";
      defparam ii2257.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2258 ( .DX(nn2258), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2257), .F2(dummy_abc_1389_), .F3(dummy_abc_1390_) );
      defparam ii2258.CONFIG_DATA = 16'h9999;
      defparam ii2258.PLACE_LOCATION = "NONE";
      defparam ii2258.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2259 ( .DX(nn2259), .F0(nn2207), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_6|SUM_net ), .F3(dummy_abc_1391_) );
      defparam ii2259.CONFIG_DATA = 16'hB8B8;
      defparam ii2259.PLACE_LOCATION = "NONE";
      defparam ii2259.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2260 ( .DX(nn2260), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2259), .F2(dummy_abc_1392_), .F3(dummy_abc_1393_) );
      defparam ii2260.CONFIG_DATA = 16'h9999;
      defparam ii2260.PLACE_LOCATION = "NONE";
      defparam ii2260.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2261 ( .DX(nn2261), .F0(nn2208), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_7|SUM_net ), .F3(dummy_abc_1394_) );
      defparam ii2261.CONFIG_DATA = 16'hB8B8;
      defparam ii2261.PLACE_LOCATION = "NONE";
      defparam ii2261.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2262 ( .DX(nn2262), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2261), .F2(dummy_abc_1395_), .F3(dummy_abc_1396_) );
      defparam ii2262.CONFIG_DATA = 16'h9999;
      defparam ii2262.PLACE_LOCATION = "NONE";
      defparam ii2262.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2263 ( .DX(nn2263), .F0(nn2209), .F1(dummy_698_), .F2(\coefcal1_divide_inst2_u110_XORCI_8|SUM_net ), .F3(dummy_abc_1397_) );
      defparam ii2263.CONFIG_DATA = 16'hB8B8;
      defparam ii2263.PLACE_LOCATION = "NONE";
      defparam ii2263.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2264 ( .DX(nn2264), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2263), .F2(dummy_abc_1398_), .F3(dummy_abc_1399_) );
      defparam ii2264.CONFIG_DATA = 16'h9999;
      defparam ii2264.PLACE_LOCATION = "NONE";
      defparam ii2264.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2265 ( .DX(nn2265), .F0(dummy_679_), .F1(\coefcal1_divide_inst2_u109_XORCI_8|SUM_net ), .F2(dummy_abc_1400_), .F3(dummy_abc_1401_) );
      defparam ii2265.CONFIG_DATA = 16'h1111;
      defparam ii2265.PLACE_LOCATION = "NONE";
      defparam ii2265.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2266 ( .DX(nn2266), .F0(nn2081), .F1(nn2265), .F2(dummy_698_), .F3(\coefcal1_divide_inst2_u110_XORCI_9|SUM_net ) );
      defparam ii2266.CONFIG_DATA = 16'h2A20;
      defparam ii2266.PLACE_LOCATION = "NONE";
      defparam ii2266.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2267 ( .DX(nn2267), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2266), .F2(dummy_abc_1402_), .F3(dummy_abc_1403_) );
      defparam ii2267.CONFIG_DATA = 16'h9999;
      defparam ii2267.PLACE_LOCATION = "NONE";
      defparam ii2267.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2268 ( .DX(nn2268), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1404_), .F2(dummy_abc_1405_), .F3(dummy_abc_1406_) );
      defparam ii2268.CONFIG_DATA = 16'h5555;
      defparam ii2268.PLACE_LOCATION = "NONE";
      defparam ii2268.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2269 ( .DX(nn2269), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1407_), .F2(dummy_abc_1408_), .F3(dummy_abc_1409_) );
      defparam ii2269.CONFIG_DATA = 16'h5555;
      defparam ii2269.PLACE_LOCATION = "NONE";
      defparam ii2269.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2270 ( .DX(nn2270), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1410_), .F2(dummy_abc_1411_), .F3(dummy_abc_1412_) );
      defparam ii2270.CONFIG_DATA = 16'h5555;
      defparam ii2270.PLACE_LOCATION = "NONE";
      defparam ii2270.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2271 ( .DX(nn2271), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1413_), .F2(dummy_abc_1414_), .F3(dummy_abc_1415_) );
      defparam ii2271.CONFIG_DATA = 16'h5555;
      defparam ii2271.PLACE_LOCATION = "NONE";
      defparam ii2271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2272 ( .DX(nn2272), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1416_), .F2(dummy_abc_1417_), .F3(dummy_abc_1418_) );
      defparam ii2272.CONFIG_DATA = 16'h5555;
      defparam ii2272.PLACE_LOCATION = "NONE";
      defparam ii2272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2273 ( .DX(nn2273), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1419_), .F2(dummy_abc_1420_), .F3(dummy_abc_1421_) );
      defparam ii2273.CONFIG_DATA = 16'h5555;
      defparam ii2273.PLACE_LOCATION = "NONE";
      defparam ii2273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2274 ( .DX(nn2274), .F0(dummy_abc_1422_), .F1(dummy_abc_1423_), .F2(dummy_abc_1424_), .F3(dummy_abc_1425_) );
      defparam ii2274.CONFIG_DATA = 16'hFFFF;
      defparam ii2274.PLACE_LOCATION = "NONE";
      defparam ii2274.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_270_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_717_ ), 
        .DX( {nn2274, nn2273, nn2272, nn2271, nn2270, nn2269, nn2268, nn2267, 
              nn2264, nn2262, nn2260, nn2258, nn2256, nn2254, nn2252, nn2250, 
              nn2248, nn2247} ), 
        .SUM( {\coefcal1_divide_inst2_u138_XORCI_17|SUM_net , dummy_718_, 
              dummy_719_, dummy_720_, dummy_721_, dummy_722_, dummy_723_, dummy_724_, 
              dummy_725_, dummy_726_, dummy_727_, dummy_728_, dummy_729_, dummy_730_, 
              dummy_731_, dummy_732_, dummy_733_, dummy_734_} )
      );
    CS_LUT4_PRIM ii2295 ( .DX(nn2295), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_698_), .F3(dummy_abc_1426_) );
      defparam ii2295.CONFIG_DATA = 16'hA6A6;
      defparam ii2295.PLACE_LOCATION = "NONE";
      defparam ii2295.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2296 ( .DX(nn2296), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1427_), .F3(dummy_abc_1428_) );
      defparam ii2296.CONFIG_DATA = 16'h9999;
      defparam ii2296.PLACE_LOCATION = "NONE";
      defparam ii2296.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2297 ( .DX(nn2297), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_698_) );
      defparam ii2297.CONFIG_DATA = 16'hA569;
      defparam ii2297.PLACE_LOCATION = "NONE";
      defparam ii2297.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2298 ( .DX(nn2298), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2249), .F2(dummy_abc_1429_), .F3(dummy_abc_1430_) );
      defparam ii2298.CONFIG_DATA = 16'h9999;
      defparam ii2298.PLACE_LOCATION = "NONE";
      defparam ii2298.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2299 ( .DX(nn2299), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2251), .F2(dummy_abc_1431_), .F3(dummy_abc_1432_) );
      defparam ii2299.CONFIG_DATA = 16'h9999;
      defparam ii2299.PLACE_LOCATION = "NONE";
      defparam ii2299.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2300 ( .DX(nn2300), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2253), .F2(dummy_abc_1433_), .F3(dummy_abc_1434_) );
      defparam ii2300.CONFIG_DATA = 16'h9999;
      defparam ii2300.PLACE_LOCATION = "NONE";
      defparam ii2300.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2301 ( .DX(nn2301), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2255), .F2(dummy_abc_1435_), .F3(dummy_abc_1436_) );
      defparam ii2301.CONFIG_DATA = 16'h9999;
      defparam ii2301.PLACE_LOCATION = "NONE";
      defparam ii2301.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2302 ( .DX(nn2302), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2257), .F2(dummy_abc_1437_), .F3(dummy_abc_1438_) );
      defparam ii2302.CONFIG_DATA = 16'h9999;
      defparam ii2302.PLACE_LOCATION = "NONE";
      defparam ii2302.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2303 ( .DX(nn2303), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2259), .F2(dummy_abc_1439_), .F3(dummy_abc_1440_) );
      defparam ii2303.CONFIG_DATA = 16'h9999;
      defparam ii2303.PLACE_LOCATION = "NONE";
      defparam ii2303.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2304 ( .DX(nn2304), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2261), .F2(dummy_abc_1441_), .F3(dummy_abc_1442_) );
      defparam ii2304.CONFIG_DATA = 16'h9999;
      defparam ii2304.PLACE_LOCATION = "NONE";
      defparam ii2304.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2305 ( .DX(nn2305), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2263), .F2(dummy_abc_1443_), .F3(dummy_abc_1444_) );
      defparam ii2305.CONFIG_DATA = 16'h9999;
      defparam ii2305.PLACE_LOCATION = "NONE";
      defparam ii2305.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2306 ( .DX(nn2306), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2266), .F2(dummy_abc_1445_), .F3(dummy_abc_1446_) );
      defparam ii2306.CONFIG_DATA = 16'h9999;
      defparam ii2306.PLACE_LOCATION = "NONE";
      defparam ii2306.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2307 ( .DX(nn2307), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(dummy_abc_1447_), .F2(dummy_abc_1448_), .F3(dummy_abc_1449_) );
      defparam ii2307.CONFIG_DATA = 16'h5555;
      defparam ii2307.PLACE_LOCATION = "NONE";
      defparam ii2307.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2308 ( .DX(nn2308), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1450_), .F2(dummy_abc_1451_), .F3(dummy_abc_1452_) );
      defparam ii2308.CONFIG_DATA = 16'h5555;
      defparam ii2308.PLACE_LOCATION = "NONE";
      defparam ii2308.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2309 ( .DX(nn2309), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1453_), .F2(dummy_abc_1454_), .F3(dummy_abc_1455_) );
      defparam ii2309.CONFIG_DATA = 16'h5555;
      defparam ii2309.PLACE_LOCATION = "NONE";
      defparam ii2309.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2310 ( .DX(nn2310), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1456_), .F2(dummy_abc_1457_), .F3(dummy_abc_1458_) );
      defparam ii2310.CONFIG_DATA = 16'h5555;
      defparam ii2310.PLACE_LOCATION = "NONE";
      defparam ii2310.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2311 ( .DX(nn2311), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1459_), .F2(dummy_abc_1460_), .F3(dummy_abc_1461_) );
      defparam ii2311.CONFIG_DATA = 16'h5555;
      defparam ii2311.PLACE_LOCATION = "NONE";
      defparam ii2311.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2312 ( .DX(nn2312), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1462_), .F2(dummy_abc_1463_), .F3(dummy_abc_1464_) );
      defparam ii2312.CONFIG_DATA = 16'h5555;
      defparam ii2312.PLACE_LOCATION = "NONE";
      defparam ii2312.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_254_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn2266, nn2263, nn2261, nn2259, nn2257, nn2255, nn2253, 
              nn2251, nn2249, nn2295, \coefcal1_yDividend__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_189_ ), 
        .DX( {nn2312, nn2311, nn2310, nn2309, nn2308, nn2307, nn2306, nn2305, 
              nn2304, nn2303, nn2302, nn2301, nn2300, nn2299, nn2298, nn2297, 
              nn2296} ), 
        .SUM( {dummy_190_, \coefcal1_divide_inst2_u111_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_14|SUM_net , \coefcal1_divide_inst2_u111_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_12|SUM_net , \coefcal1_divide_inst2_u111_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_10|SUM_net , \coefcal1_divide_inst2_u111_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_8|SUM_net , \coefcal1_divide_inst2_u111_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_6|SUM_net , \coefcal1_divide_inst2_u111_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_4|SUM_net , \coefcal1_divide_inst2_u111_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_2|SUM_net , \coefcal1_divide_inst2_u111_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2332 ( .DX(nn2332), .F0(nn2081), .F1(nn2246), .F2(dummy_717_), .F3(\coefcal1_divide_inst2_u111_XORCI_10|SUM_net ) );
      defparam ii2332.CONFIG_DATA = 16'h8A80;
      defparam ii2332.PLACE_LOCATION = "NONE";
      defparam ii2332.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2333 ( .DX(nn2333), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1465_), .F3(dummy_abc_1466_) );
      defparam ii2333.CONFIG_DATA = 16'h9999;
      defparam ii2333.PLACE_LOCATION = "NONE";
      defparam ii2333.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2334 ( .DX(nn2334), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_717_) );
      defparam ii2334.CONFIG_DATA = 16'hA569;
      defparam ii2334.PLACE_LOCATION = "NONE";
      defparam ii2334.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2335 ( .DX(nn2335), .F0(dummy_717_), .F1(nn2295), .F2(\coefcal1_divide_inst2_u111_XORCI_1|SUM_net ), .F3(dummy_abc_1467_) );
      defparam ii2335.CONFIG_DATA = 16'hD8D8;
      defparam ii2335.PLACE_LOCATION = "NONE";
      defparam ii2335.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2336 ( .DX(nn2336), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2335), .F2(dummy_abc_1468_), .F3(dummy_abc_1469_) );
      defparam ii2336.CONFIG_DATA = 16'h9999;
      defparam ii2336.PLACE_LOCATION = "NONE";
      defparam ii2336.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2337 ( .DX(nn2337), .F0(nn2249), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_2|SUM_net ), .F3(dummy_abc_1470_) );
      defparam ii2337.CONFIG_DATA = 16'hB8B8;
      defparam ii2337.PLACE_LOCATION = "NONE";
      defparam ii2337.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2338 ( .DX(nn2338), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2337), .F2(dummy_abc_1471_), .F3(dummy_abc_1472_) );
      defparam ii2338.CONFIG_DATA = 16'h9999;
      defparam ii2338.PLACE_LOCATION = "NONE";
      defparam ii2338.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2339 ( .DX(nn2339), .F0(nn2251), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_3|SUM_net ), .F3(dummy_abc_1473_) );
      defparam ii2339.CONFIG_DATA = 16'hB8B8;
      defparam ii2339.PLACE_LOCATION = "NONE";
      defparam ii2339.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2340 ( .DX(nn2340), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2339), .F2(dummy_abc_1474_), .F3(dummy_abc_1475_) );
      defparam ii2340.CONFIG_DATA = 16'h9999;
      defparam ii2340.PLACE_LOCATION = "NONE";
      defparam ii2340.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2341 ( .DX(nn2341), .F0(nn2253), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_4|SUM_net ), .F3(dummy_abc_1476_) );
      defparam ii2341.CONFIG_DATA = 16'hB8B8;
      defparam ii2341.PLACE_LOCATION = "NONE";
      defparam ii2341.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2342 ( .DX(nn2342), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2341), .F2(dummy_abc_1477_), .F3(dummy_abc_1478_) );
      defparam ii2342.CONFIG_DATA = 16'h9999;
      defparam ii2342.PLACE_LOCATION = "NONE";
      defparam ii2342.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2343 ( .DX(nn2343), .F0(nn2255), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_5|SUM_net ), .F3(dummy_abc_1479_) );
      defparam ii2343.CONFIG_DATA = 16'hB8B8;
      defparam ii2343.PLACE_LOCATION = "NONE";
      defparam ii2343.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2344 ( .DX(nn2344), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2343), .F2(dummy_abc_1480_), .F3(dummy_abc_1481_) );
      defparam ii2344.CONFIG_DATA = 16'h9999;
      defparam ii2344.PLACE_LOCATION = "NONE";
      defparam ii2344.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2345 ( .DX(nn2345), .F0(nn2257), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_6|SUM_net ), .F3(dummy_abc_1482_) );
      defparam ii2345.CONFIG_DATA = 16'hB8B8;
      defparam ii2345.PLACE_LOCATION = "NONE";
      defparam ii2345.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2346 ( .DX(nn2346), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2345), .F2(dummy_abc_1483_), .F3(dummy_abc_1484_) );
      defparam ii2346.CONFIG_DATA = 16'h9999;
      defparam ii2346.PLACE_LOCATION = "NONE";
      defparam ii2346.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2347 ( .DX(nn2347), .F0(nn2259), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_7|SUM_net ), .F3(dummy_abc_1485_) );
      defparam ii2347.CONFIG_DATA = 16'hB8B8;
      defparam ii2347.PLACE_LOCATION = "NONE";
      defparam ii2347.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2348 ( .DX(nn2348), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2347), .F2(dummy_abc_1486_), .F3(dummy_abc_1487_) );
      defparam ii2348.CONFIG_DATA = 16'h9999;
      defparam ii2348.PLACE_LOCATION = "NONE";
      defparam ii2348.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2349 ( .DX(nn2349), .F0(nn2261), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_8|SUM_net ), .F3(dummy_abc_1488_) );
      defparam ii2349.CONFIG_DATA = 16'hB8B8;
      defparam ii2349.PLACE_LOCATION = "NONE";
      defparam ii2349.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2350 ( .DX(nn2350), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2349), .F2(dummy_abc_1489_), .F3(dummy_abc_1490_) );
      defparam ii2350.CONFIG_DATA = 16'h9999;
      defparam ii2350.PLACE_LOCATION = "NONE";
      defparam ii2350.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2351 ( .DX(nn2351), .F0(nn2263), .F1(dummy_717_), .F2(\coefcal1_divide_inst2_u111_XORCI_9|SUM_net ), .F3(dummy_abc_1491_) );
      defparam ii2351.CONFIG_DATA = 16'hB8B8;
      defparam ii2351.PLACE_LOCATION = "NONE";
      defparam ii2351.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2352 ( .DX(nn2352), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2351), .F2(dummy_abc_1492_), .F3(dummy_abc_1493_) );
      defparam ii2352.CONFIG_DATA = 16'h9999;
      defparam ii2352.PLACE_LOCATION = "NONE";
      defparam ii2352.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2353 ( .DX(nn2353), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2332), .F2(dummy_abc_1494_), .F3(dummy_abc_1495_) );
      defparam ii2353.CONFIG_DATA = 16'h9999;
      defparam ii2353.PLACE_LOCATION = "NONE";
      defparam ii2353.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2354 ( .DX(nn2354), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1496_), .F2(dummy_abc_1497_), .F3(dummy_abc_1498_) );
      defparam ii2354.CONFIG_DATA = 16'h5555;
      defparam ii2354.PLACE_LOCATION = "NONE";
      defparam ii2354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2355 ( .DX(nn2355), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1499_), .F2(dummy_abc_1500_), .F3(dummy_abc_1501_) );
      defparam ii2355.CONFIG_DATA = 16'h5555;
      defparam ii2355.PLACE_LOCATION = "NONE";
      defparam ii2355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2356 ( .DX(nn2356), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1502_), .F2(dummy_abc_1503_), .F3(dummy_abc_1504_) );
      defparam ii2356.CONFIG_DATA = 16'h5555;
      defparam ii2356.PLACE_LOCATION = "NONE";
      defparam ii2356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2357 ( .DX(nn2357), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1505_), .F2(dummy_abc_1506_), .F3(dummy_abc_1507_) );
      defparam ii2357.CONFIG_DATA = 16'h5555;
      defparam ii2357.PLACE_LOCATION = "NONE";
      defparam ii2357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2358 ( .DX(nn2358), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1508_), .F2(dummy_abc_1509_), .F3(dummy_abc_1510_) );
      defparam ii2358.CONFIG_DATA = 16'h5555;
      defparam ii2358.PLACE_LOCATION = "NONE";
      defparam ii2358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2359 ( .DX(nn2359), .F0(dummy_abc_1511_), .F1(dummy_abc_1512_), .F2(dummy_abc_1513_), .F3(dummy_abc_1514_) );
      defparam ii2359.CONFIG_DATA = 16'hFFFF;
      defparam ii2359.PLACE_LOCATION = "NONE";
      defparam ii2359.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_271_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_736_ ), 
        .DX( {nn2359, nn2358, nn2357, nn2356, nn2355, nn2354, nn2353, nn2352, 
              nn2350, nn2348, nn2346, nn2344, nn2342, nn2340, nn2338, nn2336, 
              nn2334, nn2333} ), 
        .SUM( {\coefcal1_divide_inst2_u140_XORCI_17|SUM_net , dummy_737_, 
              dummy_738_, dummy_739_, dummy_740_, dummy_741_, dummy_742_, dummy_743_, 
              dummy_744_, dummy_745_, dummy_746_, dummy_747_, dummy_748_, dummy_749_, 
              dummy_750_, dummy_751_, dummy_752_, dummy_753_} )
      );
    CS_LUT4_PRIM ii2380 ( .DX(nn2380), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1515_), .F3(dummy_abc_1516_) );
      defparam ii2380.CONFIG_DATA = 16'h9999;
      defparam ii2380.PLACE_LOCATION = "NONE";
      defparam ii2380.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2381 ( .DX(nn2381), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_736_) );
      defparam ii2381.CONFIG_DATA = 16'hA569;
      defparam ii2381.PLACE_LOCATION = "NONE";
      defparam ii2381.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2382 ( .DX(nn2382), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_717_), .F3(dummy_abc_1517_) );
      defparam ii2382.CONFIG_DATA = 16'hA6A6;
      defparam ii2382.PLACE_LOCATION = "NONE";
      defparam ii2382.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2383 ( .DX(nn2383), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1518_), .F3(dummy_abc_1519_) );
      defparam ii2383.CONFIG_DATA = 16'h9999;
      defparam ii2383.PLACE_LOCATION = "NONE";
      defparam ii2383.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2384 ( .DX(nn2384), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_717_) );
      defparam ii2384.CONFIG_DATA = 16'hA569;
      defparam ii2384.PLACE_LOCATION = "NONE";
      defparam ii2384.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2385 ( .DX(nn2385), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(nn2335), .F2(dummy_abc_1520_), .F3(dummy_abc_1521_) );
      defparam ii2385.CONFIG_DATA = 16'h9999;
      defparam ii2385.PLACE_LOCATION = "NONE";
      defparam ii2385.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2386 ( .DX(nn2386), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2337), .F2(dummy_abc_1522_), .F3(dummy_abc_1523_) );
      defparam ii2386.CONFIG_DATA = 16'h9999;
      defparam ii2386.PLACE_LOCATION = "NONE";
      defparam ii2386.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2387 ( .DX(nn2387), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2339), .F2(dummy_abc_1524_), .F3(dummy_abc_1525_) );
      defparam ii2387.CONFIG_DATA = 16'h9999;
      defparam ii2387.PLACE_LOCATION = "NONE";
      defparam ii2387.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2388 ( .DX(nn2388), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2341), .F2(dummy_abc_1526_), .F3(dummy_abc_1527_) );
      defparam ii2388.CONFIG_DATA = 16'h9999;
      defparam ii2388.PLACE_LOCATION = "NONE";
      defparam ii2388.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2389 ( .DX(nn2389), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2343), .F2(dummy_abc_1528_), .F3(dummy_abc_1529_) );
      defparam ii2389.CONFIG_DATA = 16'h9999;
      defparam ii2389.PLACE_LOCATION = "NONE";
      defparam ii2389.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2390 ( .DX(nn2390), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2345), .F2(dummy_abc_1530_), .F3(dummy_abc_1531_) );
      defparam ii2390.CONFIG_DATA = 16'h9999;
      defparam ii2390.PLACE_LOCATION = "NONE";
      defparam ii2390.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2391 ( .DX(nn2391), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2347), .F2(dummy_abc_1532_), .F3(dummy_abc_1533_) );
      defparam ii2391.CONFIG_DATA = 16'h9999;
      defparam ii2391.PLACE_LOCATION = "NONE";
      defparam ii2391.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2392 ( .DX(nn2392), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2349), .F2(dummy_abc_1534_), .F3(dummy_abc_1535_) );
      defparam ii2392.CONFIG_DATA = 16'h9999;
      defparam ii2392.PLACE_LOCATION = "NONE";
      defparam ii2392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2393 ( .DX(nn2393), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2351), .F2(dummy_abc_1536_), .F3(dummy_abc_1537_) );
      defparam ii2393.CONFIG_DATA = 16'h9999;
      defparam ii2393.PLACE_LOCATION = "NONE";
      defparam ii2393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2394 ( .DX(nn2394), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2332), .F2(dummy_abc_1538_), .F3(dummy_abc_1539_) );
      defparam ii2394.CONFIG_DATA = 16'h9999;
      defparam ii2394.PLACE_LOCATION = "NONE";
      defparam ii2394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2395 ( .DX(nn2395), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_abc_1540_), .F2(dummy_abc_1541_), .F3(dummy_abc_1542_) );
      defparam ii2395.CONFIG_DATA = 16'h5555;
      defparam ii2395.PLACE_LOCATION = "NONE";
      defparam ii2395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2396 ( .DX(nn2396), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1543_), .F2(dummy_abc_1544_), .F3(dummy_abc_1545_) );
      defparam ii2396.CONFIG_DATA = 16'h5555;
      defparam ii2396.PLACE_LOCATION = "NONE";
      defparam ii2396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2397 ( .DX(nn2397), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1546_), .F2(dummy_abc_1547_), .F3(dummy_abc_1548_) );
      defparam ii2397.CONFIG_DATA = 16'h5555;
      defparam ii2397.PLACE_LOCATION = "NONE";
      defparam ii2397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2398 ( .DX(nn2398), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1549_), .F2(dummy_abc_1550_), .F3(dummy_abc_1551_) );
      defparam ii2398.CONFIG_DATA = 16'h5555;
      defparam ii2398.PLACE_LOCATION = "NONE";
      defparam ii2398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2399 ( .DX(nn2399), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1552_), .F2(dummy_abc_1553_), .F3(dummy_abc_1554_) );
      defparam ii2399.CONFIG_DATA = 16'h5555;
      defparam ii2399.PLACE_LOCATION = "NONE";
      defparam ii2399.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_255_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn2332, 
              nn2351, nn2349, nn2347, nn2345, nn2343, nn2341, nn2339, nn2337, 
              nn2335, nn2382, \coefcal1_yDividend__reg[5]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_191_ ), 
        .DX( {nn2399, nn2398, nn2397, nn2396, nn2395, nn2394, nn2393, nn2392, 
              nn2391, nn2390, nn2389, nn2388, nn2387, nn2386, nn2385, nn2384, 
              nn2383} ), 
        .SUM( {dummy_192_, \coefcal1_divide_inst2_u112_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_14|SUM_net , \coefcal1_divide_inst2_u112_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_12|SUM_net , \coefcal1_divide_inst2_u112_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_10|SUM_net , \coefcal1_divide_inst2_u112_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_8|SUM_net , \coefcal1_divide_inst2_u112_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_6|SUM_net , \coefcal1_divide_inst2_u112_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_4|SUM_net , \coefcal1_divide_inst2_u112_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_2|SUM_net , \coefcal1_divide_inst2_u112_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2419 ( .DX(nn2419), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_736_), .F2(nn2382), .F3(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ) );
      defparam ii2419.CONFIG_DATA = 16'hA695;
      defparam ii2419.PLACE_LOCATION = "NONE";
      defparam ii2419.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2420 ( .DX(nn2420), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2335), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ) );
      defparam ii2420.CONFIG_DATA = 16'h9A95;
      defparam ii2420.PLACE_LOCATION = "NONE";
      defparam ii2420.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2421 ( .DX(nn2421), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2337), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ) );
      defparam ii2421.CONFIG_DATA = 16'h9A95;
      defparam ii2421.PLACE_LOCATION = "NONE";
      defparam ii2421.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2422 ( .DX(nn2422), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2339), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ) );
      defparam ii2422.CONFIG_DATA = 16'h9A95;
      defparam ii2422.PLACE_LOCATION = "NONE";
      defparam ii2422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2423 ( .DX(nn2423), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2341), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ) );
      defparam ii2423.CONFIG_DATA = 16'h9A95;
      defparam ii2423.PLACE_LOCATION = "NONE";
      defparam ii2423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2424 ( .DX(nn2424), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2343), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ) );
      defparam ii2424.CONFIG_DATA = 16'h9A95;
      defparam ii2424.PLACE_LOCATION = "NONE";
      defparam ii2424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2425 ( .DX(nn2425), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2345), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ) );
      defparam ii2425.CONFIG_DATA = 16'h9A95;
      defparam ii2425.PLACE_LOCATION = "NONE";
      defparam ii2425.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2426 ( .DX(nn2426), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2347), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ) );
      defparam ii2426.CONFIG_DATA = 16'h9A95;
      defparam ii2426.PLACE_LOCATION = "NONE";
      defparam ii2426.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2427 ( .DX(nn2427), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2349), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ) );
      defparam ii2427.CONFIG_DATA = 16'h9A95;
      defparam ii2427.PLACE_LOCATION = "NONE";
      defparam ii2427.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2428 ( .DX(nn2428), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2351), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ) );
      defparam ii2428.CONFIG_DATA = 16'h9A95;
      defparam ii2428.PLACE_LOCATION = "NONE";
      defparam ii2428.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2429 ( .DX(nn2429), .F0(nn2332), .F1(dummy_736_), .F2(dummy_abc_1555_), .F3(dummy_abc_1556_) );
      defparam ii2429.CONFIG_DATA = 16'h8888;
      defparam ii2429.PLACE_LOCATION = "NONE";
      defparam ii2429.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2430 ( .DX(nn2430), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_11|SUM_net ), .F3(nn2429) );
      defparam ii2430.CONFIG_DATA = 16'hAA65;
      defparam ii2430.PLACE_LOCATION = "NONE";
      defparam ii2430.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2431 ( .DX(nn2431), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1557_), .F2(dummy_abc_1558_), .F3(dummy_abc_1559_) );
      defparam ii2431.CONFIG_DATA = 16'h5555;
      defparam ii2431.PLACE_LOCATION = "NONE";
      defparam ii2431.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2432 ( .DX(nn2432), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1560_), .F2(dummy_abc_1561_), .F3(dummy_abc_1562_) );
      defparam ii2432.CONFIG_DATA = 16'h5555;
      defparam ii2432.PLACE_LOCATION = "NONE";
      defparam ii2432.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2433 ( .DX(nn2433), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1563_), .F2(dummy_abc_1564_), .F3(dummy_abc_1565_) );
      defparam ii2433.CONFIG_DATA = 16'h5555;
      defparam ii2433.PLACE_LOCATION = "NONE";
      defparam ii2433.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2434 ( .DX(nn2434), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1566_), .F2(dummy_abc_1567_), .F3(dummy_abc_1568_) );
      defparam ii2434.CONFIG_DATA = 16'h5555;
      defparam ii2434.PLACE_LOCATION = "NONE";
      defparam ii2434.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2435 ( .DX(nn2435), .F0(dummy_abc_1569_), .F1(dummy_abc_1570_), .F2(dummy_abc_1571_), .F3(dummy_abc_1572_) );
      defparam ii2435.CONFIG_DATA = 16'hFFFF;
      defparam ii2435.PLACE_LOCATION = "NONE";
      defparam ii2435.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_272_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_755_ ), 
        .DX( {nn2435, nn2434, nn2433, nn2432, nn2431, nn2430, nn2428, nn2427, 
              nn2426, nn2425, nn2424, nn2423, nn2422, nn2421, nn2420, nn2419, 
              nn2381, nn2380} ), 
        .SUM( {\coefcal1_divide_inst2_u142_XORCI_17|SUM_net , dummy_756_, 
              dummy_757_, dummy_758_, dummy_759_, dummy_760_, dummy_761_, dummy_762_, 
              dummy_763_, dummy_764_, dummy_765_, dummy_766_, dummy_767_, dummy_768_, 
              dummy_769_, dummy_770_, dummy_771_, dummy_772_} )
      );
    CS_LUT4_PRIM ii2456 ( .DX(nn2456), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_736_), .F3(dummy_abc_1573_) );
      defparam ii2456.CONFIG_DATA = 16'hA6A6;
      defparam ii2456.PLACE_LOCATION = "NONE";
      defparam ii2456.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2457 ( .DX(nn2457), .F0(dummy_736_), .F1(nn2382), .F2(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ), .F3(dummy_abc_1574_) );
      defparam ii2457.CONFIG_DATA = 16'hD8D8;
      defparam ii2457.PLACE_LOCATION = "NONE";
      defparam ii2457.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2458 ( .DX(nn2458), .F0(nn2335), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ), .F3(dummy_abc_1575_) );
      defparam ii2458.CONFIG_DATA = 16'hB8B8;
      defparam ii2458.PLACE_LOCATION = "NONE";
      defparam ii2458.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2459 ( .DX(nn2459), .F0(nn2337), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ), .F3(dummy_abc_1576_) );
      defparam ii2459.CONFIG_DATA = 16'hB8B8;
      defparam ii2459.PLACE_LOCATION = "NONE";
      defparam ii2459.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2460 ( .DX(nn2460), .F0(nn2339), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ), .F3(dummy_abc_1577_) );
      defparam ii2460.CONFIG_DATA = 16'hB8B8;
      defparam ii2460.PLACE_LOCATION = "NONE";
      defparam ii2460.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2461 ( .DX(nn2461), .F0(nn2341), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ), .F3(dummy_abc_1578_) );
      defparam ii2461.CONFIG_DATA = 16'hB8B8;
      defparam ii2461.PLACE_LOCATION = "NONE";
      defparam ii2461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2462 ( .DX(nn2462), .F0(nn2343), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ), .F3(dummy_abc_1579_) );
      defparam ii2462.CONFIG_DATA = 16'hB8B8;
      defparam ii2462.PLACE_LOCATION = "NONE";
      defparam ii2462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2463 ( .DX(nn2463), .F0(nn2345), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ), .F3(dummy_abc_1580_) );
      defparam ii2463.CONFIG_DATA = 16'hB8B8;
      defparam ii2463.PLACE_LOCATION = "NONE";
      defparam ii2463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2464 ( .DX(nn2464), .F0(nn2347), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ), .F3(dummy_abc_1581_) );
      defparam ii2464.CONFIG_DATA = 16'hB8B8;
      defparam ii2464.PLACE_LOCATION = "NONE";
      defparam ii2464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2465 ( .DX(nn2465), .F0(nn2349), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ), .F3(dummy_abc_1582_) );
      defparam ii2465.CONFIG_DATA = 16'hB8B8;
      defparam ii2465.PLACE_LOCATION = "NONE";
      defparam ii2465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2466 ( .DX(nn2466), .F0(nn2351), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ), .F3(dummy_abc_1583_) );
      defparam ii2466.CONFIG_DATA = 16'hB8B8;
      defparam ii2466.PLACE_LOCATION = "NONE";
      defparam ii2466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2467 ( .DX(nn2467), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1584_), .F3(dummy_abc_1585_) );
      defparam ii2467.CONFIG_DATA = 16'h9999;
      defparam ii2467.PLACE_LOCATION = "NONE";
      defparam ii2467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2468 ( .DX(nn2468), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_736_) );
      defparam ii2468.CONFIG_DATA = 16'hA569;
      defparam ii2468.PLACE_LOCATION = "NONE";
      defparam ii2468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2469 ( .DX(nn2469), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_736_), .F2(nn2382), .F3(\coefcal1_divide_inst2_u112_XORCI_1|SUM_net ) );
      defparam ii2469.CONFIG_DATA = 16'hA695;
      defparam ii2469.PLACE_LOCATION = "NONE";
      defparam ii2469.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2470 ( .DX(nn2470), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2335), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_2|SUM_net ) );
      defparam ii2470.CONFIG_DATA = 16'h9A95;
      defparam ii2470.PLACE_LOCATION = "NONE";
      defparam ii2470.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2471 ( .DX(nn2471), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2337), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_3|SUM_net ) );
      defparam ii2471.CONFIG_DATA = 16'h9A95;
      defparam ii2471.PLACE_LOCATION = "NONE";
      defparam ii2471.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2472 ( .DX(nn2472), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2339), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_4|SUM_net ) );
      defparam ii2472.CONFIG_DATA = 16'h9A95;
      defparam ii2472.PLACE_LOCATION = "NONE";
      defparam ii2472.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2473 ( .DX(nn2473), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2341), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_5|SUM_net ) );
      defparam ii2473.CONFIG_DATA = 16'h9A95;
      defparam ii2473.PLACE_LOCATION = "NONE";
      defparam ii2473.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2474 ( .DX(nn2474), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2343), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_6|SUM_net ) );
      defparam ii2474.CONFIG_DATA = 16'h9A95;
      defparam ii2474.PLACE_LOCATION = "NONE";
      defparam ii2474.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2475 ( .DX(nn2475), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2345), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_7|SUM_net ) );
      defparam ii2475.CONFIG_DATA = 16'h9A95;
      defparam ii2475.PLACE_LOCATION = "NONE";
      defparam ii2475.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2476 ( .DX(nn2476), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2347), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_8|SUM_net ) );
      defparam ii2476.CONFIG_DATA = 16'h9A95;
      defparam ii2476.PLACE_LOCATION = "NONE";
      defparam ii2476.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2477 ( .DX(nn2477), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2349), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_9|SUM_net ) );
      defparam ii2477.CONFIG_DATA = 16'h9A95;
      defparam ii2477.PLACE_LOCATION = "NONE";
      defparam ii2477.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2478 ( .DX(nn2478), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2351), .F2(dummy_736_), .F3(\coefcal1_divide_inst2_u112_XORCI_10|SUM_net ) );
      defparam ii2478.CONFIG_DATA = 16'h9A95;
      defparam ii2478.PLACE_LOCATION = "NONE";
      defparam ii2478.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2479 ( .DX(nn2479), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(dummy_736_), .F2(\coefcal1_divide_inst2_u112_XORCI_11|SUM_net ), .F3(nn2429) );
      defparam ii2479.CONFIG_DATA = 16'hAA65;
      defparam ii2479.PLACE_LOCATION = "NONE";
      defparam ii2479.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2480 ( .DX(nn2480), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(dummy_abc_1586_), .F2(dummy_abc_1587_), .F3(dummy_abc_1588_) );
      defparam ii2480.CONFIG_DATA = 16'h5555;
      defparam ii2480.PLACE_LOCATION = "NONE";
      defparam ii2480.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2481 ( .DX(nn2481), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1589_), .F2(dummy_abc_1590_), .F3(dummy_abc_1591_) );
      defparam ii2481.CONFIG_DATA = 16'h5555;
      defparam ii2481.PLACE_LOCATION = "NONE";
      defparam ii2481.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2482 ( .DX(nn2482), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1592_), .F2(dummy_abc_1593_), .F3(dummy_abc_1594_) );
      defparam ii2482.CONFIG_DATA = 16'h5555;
      defparam ii2482.PLACE_LOCATION = "NONE";
      defparam ii2482.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2483 ( .DX(nn2483), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1595_), .F2(dummy_abc_1596_), .F3(dummy_abc_1597_) );
      defparam ii2483.CONFIG_DATA = 16'h5555;
      defparam ii2483.PLACE_LOCATION = "NONE";
      defparam ii2483.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_256_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn2466, 
              nn2465, nn2464, nn2463, nn2462, nn2461, nn2460, nn2459, nn2458, 
              nn2457, nn2456, \coefcal1_yDividend__reg[4]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_193_ ), 
        .DX( {nn2483, nn2482, nn2481, nn2480, nn2479, nn2478, nn2477, nn2476, 
              nn2475, nn2474, nn2473, nn2472, nn2471, nn2470, nn2469, nn2468, 
              nn2467} ), 
        .SUM( {dummy_194_, \coefcal1_divide_inst2_u113_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_14|SUM_net , \coefcal1_divide_inst2_u113_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_12|SUM_net , \coefcal1_divide_inst2_u113_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_10|SUM_net , \coefcal1_divide_inst2_u113_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_8|SUM_net , \coefcal1_divide_inst2_u113_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_6|SUM_net , \coefcal1_divide_inst2_u113_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_4|SUM_net , \coefcal1_divide_inst2_u113_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_2|SUM_net , \coefcal1_divide_inst2_u113_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u113_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2503 ( .DX(nn2503), .F0(nn2332), .F1(dummy_736_), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2503.CONFIG_DATA = 16'h8F80;
      defparam ii2503.PLACE_LOCATION = "NONE";
      defparam ii2503.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2504 ( .DX(nn2504), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1598_), .F3(dummy_abc_1599_) );
      defparam ii2504.CONFIG_DATA = 16'h9999;
      defparam ii2504.PLACE_LOCATION = "NONE";
      defparam ii2504.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2505 ( .DX(nn2505), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_755_) );
      defparam ii2505.CONFIG_DATA = 16'hA569;
      defparam ii2505.PLACE_LOCATION = "NONE";
      defparam ii2505.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2506 ( .DX(nn2506), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_755_), .F2(nn2456), .F3(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ) );
      defparam ii2506.CONFIG_DATA = 16'hA695;
      defparam ii2506.PLACE_LOCATION = "NONE";
      defparam ii2506.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2507 ( .DX(nn2507), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2457), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ) );
      defparam ii2507.CONFIG_DATA = 16'h9A95;
      defparam ii2507.PLACE_LOCATION = "NONE";
      defparam ii2507.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2508 ( .DX(nn2508), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2458), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ) );
      defparam ii2508.CONFIG_DATA = 16'h9A95;
      defparam ii2508.PLACE_LOCATION = "NONE";
      defparam ii2508.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2509 ( .DX(nn2509), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2459), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ) );
      defparam ii2509.CONFIG_DATA = 16'h9A95;
      defparam ii2509.PLACE_LOCATION = "NONE";
      defparam ii2509.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2510 ( .DX(nn2510), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2460), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ) );
      defparam ii2510.CONFIG_DATA = 16'h9A95;
      defparam ii2510.PLACE_LOCATION = "NONE";
      defparam ii2510.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2511 ( .DX(nn2511), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2461), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ) );
      defparam ii2511.CONFIG_DATA = 16'h9A95;
      defparam ii2511.PLACE_LOCATION = "NONE";
      defparam ii2511.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2512 ( .DX(nn2512), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2462), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ) );
      defparam ii2512.CONFIG_DATA = 16'h9A95;
      defparam ii2512.PLACE_LOCATION = "NONE";
      defparam ii2512.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2513 ( .DX(nn2513), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2463), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ) );
      defparam ii2513.CONFIG_DATA = 16'h9A95;
      defparam ii2513.PLACE_LOCATION = "NONE";
      defparam ii2513.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2514 ( .DX(nn2514), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2464), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ) );
      defparam ii2514.CONFIG_DATA = 16'h9A95;
      defparam ii2514.PLACE_LOCATION = "NONE";
      defparam ii2514.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2515 ( .DX(nn2515), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2465), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ) );
      defparam ii2515.CONFIG_DATA = 16'h9A95;
      defparam ii2515.PLACE_LOCATION = "NONE";
      defparam ii2515.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2516 ( .DX(nn2516), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2466), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ) );
      defparam ii2516.CONFIG_DATA = 16'h9A95;
      defparam ii2516.PLACE_LOCATION = "NONE";
      defparam ii2516.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2517 ( .DX(nn2517), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2429), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2517.CONFIG_DATA = 16'h9095;
      defparam ii2517.PLACE_LOCATION = "NONE";
      defparam ii2517.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2518 ( .DX(nn2518), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1600_), .F2(dummy_abc_1601_), .F3(dummy_abc_1602_) );
      defparam ii2518.CONFIG_DATA = 16'h5555;
      defparam ii2518.PLACE_LOCATION = "NONE";
      defparam ii2518.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2519 ( .DX(nn2519), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1603_), .F2(dummy_abc_1604_), .F3(dummy_abc_1605_) );
      defparam ii2519.CONFIG_DATA = 16'h5555;
      defparam ii2519.PLACE_LOCATION = "NONE";
      defparam ii2519.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2520 ( .DX(nn2520), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1606_), .F2(dummy_abc_1607_), .F3(dummy_abc_1608_) );
      defparam ii2520.CONFIG_DATA = 16'h5555;
      defparam ii2520.PLACE_LOCATION = "NONE";
      defparam ii2520.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2521 ( .DX(nn2521), .F0(dummy_abc_1609_), .F1(dummy_abc_1610_), .F2(dummy_abc_1611_), .F3(dummy_abc_1612_) );
      defparam ii2521.CONFIG_DATA = 16'hFFFF;
      defparam ii2521.PLACE_LOCATION = "NONE";
      defparam ii2521.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_273_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_774_ ), 
        .DX( {nn2521, nn2520, nn2519, nn2518, nn2517, nn2516, nn2515, nn2514, 
              nn2513, nn2512, nn2511, nn2510, nn2509, nn2508, nn2507, nn2506, 
              nn2505, nn2504} ), 
        .SUM( {\coefcal1_divide_inst2_u144_XORCI_17|SUM_net , dummy_775_, 
              dummy_776_, dummy_777_, dummy_778_, dummy_779_, dummy_780_, dummy_781_, 
              dummy_782_, dummy_783_, dummy_784_, dummy_785_, dummy_786_, dummy_787_, 
              dummy_788_, dummy_789_, dummy_790_, dummy_791_} )
      );
    CS_LUT4_PRIM ii2542 ( .DX(nn2542), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_755_), .F3(dummy_abc_1613_) );
      defparam ii2542.CONFIG_DATA = 16'hA6A6;
      defparam ii2542.PLACE_LOCATION = "NONE";
      defparam ii2542.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2543 ( .DX(nn2543), .F0(dummy_755_), .F1(nn2456), .F2(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ), .F3(dummy_abc_1614_) );
      defparam ii2543.CONFIG_DATA = 16'hD8D8;
      defparam ii2543.PLACE_LOCATION = "NONE";
      defparam ii2543.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2544 ( .DX(nn2544), .F0(nn2457), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ), .F3(dummy_abc_1615_) );
      defparam ii2544.CONFIG_DATA = 16'hB8B8;
      defparam ii2544.PLACE_LOCATION = "NONE";
      defparam ii2544.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2545 ( .DX(nn2545), .F0(nn2458), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ), .F3(dummy_abc_1616_) );
      defparam ii2545.CONFIG_DATA = 16'hB8B8;
      defparam ii2545.PLACE_LOCATION = "NONE";
      defparam ii2545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2546 ( .DX(nn2546), .F0(nn2459), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ), .F3(dummy_abc_1617_) );
      defparam ii2546.CONFIG_DATA = 16'hB8B8;
      defparam ii2546.PLACE_LOCATION = "NONE";
      defparam ii2546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2547 ( .DX(nn2547), .F0(nn2460), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ), .F3(dummy_abc_1618_) );
      defparam ii2547.CONFIG_DATA = 16'hB8B8;
      defparam ii2547.PLACE_LOCATION = "NONE";
      defparam ii2547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2548 ( .DX(nn2548), .F0(nn2461), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ), .F3(dummy_abc_1619_) );
      defparam ii2548.CONFIG_DATA = 16'hB8B8;
      defparam ii2548.PLACE_LOCATION = "NONE";
      defparam ii2548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2549 ( .DX(nn2549), .F0(nn2462), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ), .F3(dummy_abc_1620_) );
      defparam ii2549.CONFIG_DATA = 16'hB8B8;
      defparam ii2549.PLACE_LOCATION = "NONE";
      defparam ii2549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2550 ( .DX(nn2550), .F0(nn2463), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ), .F3(dummy_abc_1621_) );
      defparam ii2550.CONFIG_DATA = 16'hB8B8;
      defparam ii2550.PLACE_LOCATION = "NONE";
      defparam ii2550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2551 ( .DX(nn2551), .F0(nn2464), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ), .F3(dummy_abc_1622_) );
      defparam ii2551.CONFIG_DATA = 16'hB8B8;
      defparam ii2551.PLACE_LOCATION = "NONE";
      defparam ii2551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2552 ( .DX(nn2552), .F0(nn2465), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ), .F3(dummy_abc_1623_) );
      defparam ii2552.CONFIG_DATA = 16'hB8B8;
      defparam ii2552.PLACE_LOCATION = "NONE";
      defparam ii2552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2553 ( .DX(nn2553), .F0(nn2466), .F1(dummy_755_), .F2(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ), .F3(dummy_abc_1624_) );
      defparam ii2553.CONFIG_DATA = 16'hB8B8;
      defparam ii2553.PLACE_LOCATION = "NONE";
      defparam ii2553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2554 ( .DX(nn2554), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1625_), .F3(dummy_abc_1626_) );
      defparam ii2554.CONFIG_DATA = 16'h9999;
      defparam ii2554.PLACE_LOCATION = "NONE";
      defparam ii2554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2555 ( .DX(nn2555), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_755_) );
      defparam ii2555.CONFIG_DATA = 16'hA569;
      defparam ii2555.PLACE_LOCATION = "NONE";
      defparam ii2555.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2556 ( .DX(nn2556), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_755_), .F2(nn2456), .F3(\coefcal1_divide_inst2_u113_XORCI_1|SUM_net ) );
      defparam ii2556.CONFIG_DATA = 16'hA695;
      defparam ii2556.PLACE_LOCATION = "NONE";
      defparam ii2556.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2557 ( .DX(nn2557), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2457), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_2|SUM_net ) );
      defparam ii2557.CONFIG_DATA = 16'h9A95;
      defparam ii2557.PLACE_LOCATION = "NONE";
      defparam ii2557.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2558 ( .DX(nn2558), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2458), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_3|SUM_net ) );
      defparam ii2558.CONFIG_DATA = 16'h9A95;
      defparam ii2558.PLACE_LOCATION = "NONE";
      defparam ii2558.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2559 ( .DX(nn2559), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2459), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_4|SUM_net ) );
      defparam ii2559.CONFIG_DATA = 16'h9A95;
      defparam ii2559.PLACE_LOCATION = "NONE";
      defparam ii2559.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2560 ( .DX(nn2560), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2460), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_5|SUM_net ) );
      defparam ii2560.CONFIG_DATA = 16'h9A95;
      defparam ii2560.PLACE_LOCATION = "NONE";
      defparam ii2560.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2561 ( .DX(nn2561), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2461), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_6|SUM_net ) );
      defparam ii2561.CONFIG_DATA = 16'h9A95;
      defparam ii2561.PLACE_LOCATION = "NONE";
      defparam ii2561.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2562 ( .DX(nn2562), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2462), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_7|SUM_net ) );
      defparam ii2562.CONFIG_DATA = 16'h9A95;
      defparam ii2562.PLACE_LOCATION = "NONE";
      defparam ii2562.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2563 ( .DX(nn2563), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2463), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_8|SUM_net ) );
      defparam ii2563.CONFIG_DATA = 16'h9A95;
      defparam ii2563.PLACE_LOCATION = "NONE";
      defparam ii2563.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2564 ( .DX(nn2564), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2464), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_9|SUM_net ) );
      defparam ii2564.CONFIG_DATA = 16'h9A95;
      defparam ii2564.PLACE_LOCATION = "NONE";
      defparam ii2564.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2565 ( .DX(nn2565), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2465), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_10|SUM_net ) );
      defparam ii2565.CONFIG_DATA = 16'h9A95;
      defparam ii2565.PLACE_LOCATION = "NONE";
      defparam ii2565.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2566 ( .DX(nn2566), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2466), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_11|SUM_net ) );
      defparam ii2566.CONFIG_DATA = 16'h9A95;
      defparam ii2566.PLACE_LOCATION = "NONE";
      defparam ii2566.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2567 ( .DX(nn2567), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2429), .F2(dummy_755_), .F3(\coefcal1_divide_inst2_u113_XORCI_12|SUM_net ) );
      defparam ii2567.CONFIG_DATA = 16'h9095;
      defparam ii2567.PLACE_LOCATION = "NONE";
      defparam ii2567.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2568 ( .DX(nn2568), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(dummy_abc_1627_), .F2(dummy_abc_1628_), .F3(dummy_abc_1629_) );
      defparam ii2568.CONFIG_DATA = 16'h5555;
      defparam ii2568.PLACE_LOCATION = "NONE";
      defparam ii2568.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2569 ( .DX(nn2569), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1630_), .F2(dummy_abc_1631_), .F3(dummy_abc_1632_) );
      defparam ii2569.CONFIG_DATA = 16'h5555;
      defparam ii2569.PLACE_LOCATION = "NONE";
      defparam ii2569.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2570 ( .DX(nn2570), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1633_), .F2(dummy_abc_1634_), .F3(dummy_abc_1635_) );
      defparam ii2570.CONFIG_DATA = 16'h5555;
      defparam ii2570.PLACE_LOCATION = "NONE";
      defparam ii2570.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_257_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn2503, nn2553, nn2552, nn2551, nn2550, nn2549, nn2548, 
              nn2547, nn2546, nn2545, nn2544, nn2543, nn2542, 
              \coefcal1_yDividend__reg[3]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_195_ ), 
        .DX( {nn2570, nn2569, nn2568, nn2567, nn2566, nn2565, nn2564, nn2563, 
              nn2562, nn2561, nn2560, nn2559, nn2558, nn2557, nn2556, nn2555, 
              nn2554} ), 
        .SUM( {dummy_196_, \coefcal1_divide_inst2_u114_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_14|SUM_net , \coefcal1_divide_inst2_u114_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_12|SUM_net , \coefcal1_divide_inst2_u114_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_10|SUM_net , \coefcal1_divide_inst2_u114_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_8|SUM_net , \coefcal1_divide_inst2_u114_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_6|SUM_net , \coefcal1_divide_inst2_u114_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_4|SUM_net , \coefcal1_divide_inst2_u114_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_2|SUM_net , \coefcal1_divide_inst2_u114_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u114_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2590 ( .DX(nn2590), .F0(dummy_774_), .F1(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ), .F2(dummy_abc_1636_), .F3(dummy_abc_1637_) );
      defparam ii2590.CONFIG_DATA = 16'h1111;
      defparam ii2590.PLACE_LOCATION = "NONE";
      defparam ii2590.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2591 ( .DX(nn2591), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1638_), .F3(dummy_abc_1639_) );
      defparam ii2591.CONFIG_DATA = 16'h9999;
      defparam ii2591.PLACE_LOCATION = "NONE";
      defparam ii2591.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2592 ( .DX(nn2592), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_774_) );
      defparam ii2592.CONFIG_DATA = 16'hA569;
      defparam ii2592.PLACE_LOCATION = "NONE";
      defparam ii2592.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2593 ( .DX(nn2593), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_774_), .F2(nn2542), .F3(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ) );
      defparam ii2593.CONFIG_DATA = 16'hA695;
      defparam ii2593.PLACE_LOCATION = "NONE";
      defparam ii2593.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2594 ( .DX(nn2594), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2543), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ) );
      defparam ii2594.CONFIG_DATA = 16'h9A95;
      defparam ii2594.PLACE_LOCATION = "NONE";
      defparam ii2594.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2595 ( .DX(nn2595), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2544), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ) );
      defparam ii2595.CONFIG_DATA = 16'h9A95;
      defparam ii2595.PLACE_LOCATION = "NONE";
      defparam ii2595.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2596 ( .DX(nn2596), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2545), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ) );
      defparam ii2596.CONFIG_DATA = 16'h9A95;
      defparam ii2596.PLACE_LOCATION = "NONE";
      defparam ii2596.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2597 ( .DX(nn2597), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2546), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ) );
      defparam ii2597.CONFIG_DATA = 16'h9A95;
      defparam ii2597.PLACE_LOCATION = "NONE";
      defparam ii2597.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2598 ( .DX(nn2598), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2547), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ) );
      defparam ii2598.CONFIG_DATA = 16'h9A95;
      defparam ii2598.PLACE_LOCATION = "NONE";
      defparam ii2598.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2599 ( .DX(nn2599), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2548), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ) );
      defparam ii2599.CONFIG_DATA = 16'h9A95;
      defparam ii2599.PLACE_LOCATION = "NONE";
      defparam ii2599.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2600 ( .DX(nn2600), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2549), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ) );
      defparam ii2600.CONFIG_DATA = 16'h9A95;
      defparam ii2600.PLACE_LOCATION = "NONE";
      defparam ii2600.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2601 ( .DX(nn2601), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2550), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ) );
      defparam ii2601.CONFIG_DATA = 16'h9A95;
      defparam ii2601.PLACE_LOCATION = "NONE";
      defparam ii2601.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2602 ( .DX(nn2602), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2551), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ) );
      defparam ii2602.CONFIG_DATA = 16'h9A95;
      defparam ii2602.PLACE_LOCATION = "NONE";
      defparam ii2602.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2603 ( .DX(nn2603), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2552), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ) );
      defparam ii2603.CONFIG_DATA = 16'h9A95;
      defparam ii2603.PLACE_LOCATION = "NONE";
      defparam ii2603.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2604 ( .DX(nn2604), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2553), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ) );
      defparam ii2604.CONFIG_DATA = 16'h9A95;
      defparam ii2604.PLACE_LOCATION = "NONE";
      defparam ii2604.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2605 ( .DX(nn2605), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2503), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ) );
      defparam ii2605.CONFIG_DATA = 16'h9995;
      defparam ii2605.PLACE_LOCATION = "NONE";
      defparam ii2605.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2606 ( .DX(nn2606), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1640_), .F2(dummy_abc_1641_), .F3(dummy_abc_1642_) );
      defparam ii2606.CONFIG_DATA = 16'h5555;
      defparam ii2606.PLACE_LOCATION = "NONE";
      defparam ii2606.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2607 ( .DX(nn2607), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1643_), .F2(dummy_abc_1644_), .F3(dummy_abc_1645_) );
      defparam ii2607.CONFIG_DATA = 16'h5555;
      defparam ii2607.PLACE_LOCATION = "NONE";
      defparam ii2607.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2608 ( .DX(nn2608), .F0(dummy_abc_1646_), .F1(dummy_abc_1647_), .F2(dummy_abc_1648_), .F3(dummy_abc_1649_) );
      defparam ii2608.CONFIG_DATA = 16'hFFFF;
      defparam ii2608.PLACE_LOCATION = "NONE";
      defparam ii2608.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_274_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_793_ ), 
        .DX( {nn2608, nn2607, nn2606, nn2605, nn2604, nn2603, nn2602, nn2601, 
              nn2600, nn2599, nn2598, nn2597, nn2596, nn2595, nn2594, nn2593, 
              nn2592, nn2591} ), 
        .SUM( {\coefcal1_divide_inst2_u146_XORCI_17|SUM_net , dummy_794_, 
              dummy_795_, dummy_796_, dummy_797_, dummy_798_, dummy_799_, dummy_800_, 
              dummy_801_, dummy_802_, dummy_803_, dummy_804_, dummy_805_, dummy_806_, 
              dummy_807_, dummy_808_, dummy_809_, dummy_810_} )
      );
    CS_LUT4_PRIM ii2629 ( .DX(nn2629), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_774_), .F3(dummy_abc_1650_) );
      defparam ii2629.CONFIG_DATA = 16'hA6A6;
      defparam ii2629.PLACE_LOCATION = "NONE";
      defparam ii2629.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2630 ( .DX(nn2630), .F0(dummy_774_), .F1(nn2542), .F2(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ), .F3(dummy_abc_1651_) );
      defparam ii2630.CONFIG_DATA = 16'hD8D8;
      defparam ii2630.PLACE_LOCATION = "NONE";
      defparam ii2630.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2631 ( .DX(nn2631), .F0(nn2543), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ), .F3(dummy_abc_1652_) );
      defparam ii2631.CONFIG_DATA = 16'hB8B8;
      defparam ii2631.PLACE_LOCATION = "NONE";
      defparam ii2631.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2632 ( .DX(nn2632), .F0(nn2544), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ), .F3(dummy_abc_1653_) );
      defparam ii2632.CONFIG_DATA = 16'hB8B8;
      defparam ii2632.PLACE_LOCATION = "NONE";
      defparam ii2632.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2633 ( .DX(nn2633), .F0(nn2545), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ), .F3(dummy_abc_1654_) );
      defparam ii2633.CONFIG_DATA = 16'hB8B8;
      defparam ii2633.PLACE_LOCATION = "NONE";
      defparam ii2633.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2634 ( .DX(nn2634), .F0(nn2546), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ), .F3(dummy_abc_1655_) );
      defparam ii2634.CONFIG_DATA = 16'hB8B8;
      defparam ii2634.PLACE_LOCATION = "NONE";
      defparam ii2634.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2635 ( .DX(nn2635), .F0(nn2547), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ), .F3(dummy_abc_1656_) );
      defparam ii2635.CONFIG_DATA = 16'hB8B8;
      defparam ii2635.PLACE_LOCATION = "NONE";
      defparam ii2635.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2636 ( .DX(nn2636), .F0(nn2548), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ), .F3(dummy_abc_1657_) );
      defparam ii2636.CONFIG_DATA = 16'hB8B8;
      defparam ii2636.PLACE_LOCATION = "NONE";
      defparam ii2636.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2637 ( .DX(nn2637), .F0(nn2549), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ), .F3(dummy_abc_1658_) );
      defparam ii2637.CONFIG_DATA = 16'hB8B8;
      defparam ii2637.PLACE_LOCATION = "NONE";
      defparam ii2637.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2638 ( .DX(nn2638), .F0(nn2550), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ), .F3(dummy_abc_1659_) );
      defparam ii2638.CONFIG_DATA = 16'hB8B8;
      defparam ii2638.PLACE_LOCATION = "NONE";
      defparam ii2638.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2639 ( .DX(nn2639), .F0(nn2551), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ), .F3(dummy_abc_1660_) );
      defparam ii2639.CONFIG_DATA = 16'hB8B8;
      defparam ii2639.PLACE_LOCATION = "NONE";
      defparam ii2639.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2640 ( .DX(nn2640), .F0(nn2552), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ), .F3(dummy_abc_1661_) );
      defparam ii2640.CONFIG_DATA = 16'hB8B8;
      defparam ii2640.PLACE_LOCATION = "NONE";
      defparam ii2640.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2641 ( .DX(nn2641), .F0(nn2553), .F1(dummy_774_), .F2(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ), .F3(dummy_abc_1662_) );
      defparam ii2641.CONFIG_DATA = 16'hB8B8;
      defparam ii2641.PLACE_LOCATION = "NONE";
      defparam ii2641.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2642 ( .DX(nn2642), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1663_), .F3(dummy_abc_1664_) );
      defparam ii2642.CONFIG_DATA = 16'h9999;
      defparam ii2642.PLACE_LOCATION = "NONE";
      defparam ii2642.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2643 ( .DX(nn2643), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_774_) );
      defparam ii2643.CONFIG_DATA = 16'hA569;
      defparam ii2643.PLACE_LOCATION = "NONE";
      defparam ii2643.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2644 ( .DX(nn2644), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_774_), .F2(nn2542), .F3(\coefcal1_divide_inst2_u114_XORCI_1|SUM_net ) );
      defparam ii2644.CONFIG_DATA = 16'hA695;
      defparam ii2644.PLACE_LOCATION = "NONE";
      defparam ii2644.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2645 ( .DX(nn2645), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2543), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_2|SUM_net ) );
      defparam ii2645.CONFIG_DATA = 16'h9A95;
      defparam ii2645.PLACE_LOCATION = "NONE";
      defparam ii2645.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2646 ( .DX(nn2646), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2544), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_3|SUM_net ) );
      defparam ii2646.CONFIG_DATA = 16'h9A95;
      defparam ii2646.PLACE_LOCATION = "NONE";
      defparam ii2646.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2647 ( .DX(nn2647), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2545), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_4|SUM_net ) );
      defparam ii2647.CONFIG_DATA = 16'h9A95;
      defparam ii2647.PLACE_LOCATION = "NONE";
      defparam ii2647.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2648 ( .DX(nn2648), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2546), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_5|SUM_net ) );
      defparam ii2648.CONFIG_DATA = 16'h9A95;
      defparam ii2648.PLACE_LOCATION = "NONE";
      defparam ii2648.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2649 ( .DX(nn2649), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2547), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_6|SUM_net ) );
      defparam ii2649.CONFIG_DATA = 16'h9A95;
      defparam ii2649.PLACE_LOCATION = "NONE";
      defparam ii2649.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2650 ( .DX(nn2650), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2548), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_7|SUM_net ) );
      defparam ii2650.CONFIG_DATA = 16'h9A95;
      defparam ii2650.PLACE_LOCATION = "NONE";
      defparam ii2650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2651 ( .DX(nn2651), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2549), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_8|SUM_net ) );
      defparam ii2651.CONFIG_DATA = 16'h9A95;
      defparam ii2651.PLACE_LOCATION = "NONE";
      defparam ii2651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2652 ( .DX(nn2652), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2550), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_9|SUM_net ) );
      defparam ii2652.CONFIG_DATA = 16'h9A95;
      defparam ii2652.PLACE_LOCATION = "NONE";
      defparam ii2652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2653 ( .DX(nn2653), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2551), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_10|SUM_net ) );
      defparam ii2653.CONFIG_DATA = 16'h9A95;
      defparam ii2653.PLACE_LOCATION = "NONE";
      defparam ii2653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2654 ( .DX(nn2654), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2552), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_11|SUM_net ) );
      defparam ii2654.CONFIG_DATA = 16'h9A95;
      defparam ii2654.PLACE_LOCATION = "NONE";
      defparam ii2654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2655 ( .DX(nn2655), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2553), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_12|SUM_net ) );
      defparam ii2655.CONFIG_DATA = 16'h9A95;
      defparam ii2655.PLACE_LOCATION = "NONE";
      defparam ii2655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2656 ( .DX(nn2656), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2503), .F2(dummy_774_), .F3(\coefcal1_divide_inst2_u114_XORCI_13|SUM_net ) );
      defparam ii2656.CONFIG_DATA = 16'h9995;
      defparam ii2656.PLACE_LOCATION = "NONE";
      defparam ii2656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2657 ( .DX(nn2657), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(dummy_abc_1665_), .F2(dummy_abc_1666_), .F3(dummy_abc_1667_) );
      defparam ii2657.CONFIG_DATA = 16'h5555;
      defparam ii2657.PLACE_LOCATION = "NONE";
      defparam ii2657.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2658 ( .DX(nn2658), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1668_), .F2(dummy_abc_1669_), .F3(dummy_abc_1670_) );
      defparam ii2658.CONFIG_DATA = 16'h5555;
      defparam ii2658.PLACE_LOCATION = "NONE";
      defparam ii2658.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_258_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn2641, nn2640, nn2639, nn2638, nn2637, nn2636, nn2635, 
              nn2634, nn2633, nn2632, nn2631, nn2630, nn2629, 
              \coefcal1_yDividend__reg[2]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_197_ ), 
        .DX( {nn2658, nn2657, nn2656, nn2655, nn2654, nn2653, nn2652, nn2651, 
              nn2650, nn2649, nn2648, nn2647, nn2646, nn2645, nn2644, nn2643, 
              nn2642} ), 
        .SUM( {dummy_198_, \coefcal1_divide_inst2_u115_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_14|SUM_net , \coefcal1_divide_inst2_u115_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_12|SUM_net , \coefcal1_divide_inst2_u115_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_10|SUM_net , \coefcal1_divide_inst2_u115_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_8|SUM_net , \coefcal1_divide_inst2_u115_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_6|SUM_net , \coefcal1_divide_inst2_u115_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_4|SUM_net , \coefcal1_divide_inst2_u115_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_2|SUM_net , \coefcal1_divide_inst2_u115_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u115_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2678 ( .DX(nn2678), .F0(nn2503), .F1(nn2590), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_14|SUM_net ) );
      defparam ii2678.CONFIG_DATA = 16'h2A20;
      defparam ii2678.PLACE_LOCATION = "NONE";
      defparam ii2678.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2679 ( .DX(nn2679), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1671_), .F3(dummy_abc_1672_) );
      defparam ii2679.CONFIG_DATA = 16'h9999;
      defparam ii2679.PLACE_LOCATION = "NONE";
      defparam ii2679.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2680 ( .DX(nn2680), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_793_) );
      defparam ii2680.CONFIG_DATA = 16'hA569;
      defparam ii2680.PLACE_LOCATION = "NONE";
      defparam ii2680.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2681 ( .DX(nn2681), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_793_), .F2(nn2629), .F3(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ) );
      defparam ii2681.CONFIG_DATA = 16'hA695;
      defparam ii2681.PLACE_LOCATION = "NONE";
      defparam ii2681.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2682 ( .DX(nn2682), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2630), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ) );
      defparam ii2682.CONFIG_DATA = 16'h9A95;
      defparam ii2682.PLACE_LOCATION = "NONE";
      defparam ii2682.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2683 ( .DX(nn2683), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2631), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ) );
      defparam ii2683.CONFIG_DATA = 16'h9A95;
      defparam ii2683.PLACE_LOCATION = "NONE";
      defparam ii2683.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2684 ( .DX(nn2684), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2632), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ) );
      defparam ii2684.CONFIG_DATA = 16'h9A95;
      defparam ii2684.PLACE_LOCATION = "NONE";
      defparam ii2684.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2685 ( .DX(nn2685), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2633), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ) );
      defparam ii2685.CONFIG_DATA = 16'h9A95;
      defparam ii2685.PLACE_LOCATION = "NONE";
      defparam ii2685.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2686 ( .DX(nn2686), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2634), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ) );
      defparam ii2686.CONFIG_DATA = 16'h9A95;
      defparam ii2686.PLACE_LOCATION = "NONE";
      defparam ii2686.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2687 ( .DX(nn2687), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2635), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ) );
      defparam ii2687.CONFIG_DATA = 16'h9A95;
      defparam ii2687.PLACE_LOCATION = "NONE";
      defparam ii2687.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2688 ( .DX(nn2688), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2636), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ) );
      defparam ii2688.CONFIG_DATA = 16'h9A95;
      defparam ii2688.PLACE_LOCATION = "NONE";
      defparam ii2688.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2689 ( .DX(nn2689), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2637), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ) );
      defparam ii2689.CONFIG_DATA = 16'h9A95;
      defparam ii2689.PLACE_LOCATION = "NONE";
      defparam ii2689.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2690 ( .DX(nn2690), .F0(nn2638), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_10|SUM_net ), .F3(dummy_abc_1673_) );
      defparam ii2690.CONFIG_DATA = 16'hB8B8;
      defparam ii2690.PLACE_LOCATION = "NONE";
      defparam ii2690.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2691 ( .DX(nn2691), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2690), .F2(dummy_abc_1674_), .F3(dummy_abc_1675_) );
      defparam ii2691.CONFIG_DATA = 16'h9999;
      defparam ii2691.PLACE_LOCATION = "NONE";
      defparam ii2691.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2692 ( .DX(nn2692), .F0(nn2639), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_11|SUM_net ), .F3(dummy_abc_1676_) );
      defparam ii2692.CONFIG_DATA = 16'hB8B8;
      defparam ii2692.PLACE_LOCATION = "NONE";
      defparam ii2692.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2693 ( .DX(nn2693), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2692), .F2(dummy_abc_1677_), .F3(dummy_abc_1678_) );
      defparam ii2693.CONFIG_DATA = 16'h9999;
      defparam ii2693.PLACE_LOCATION = "NONE";
      defparam ii2693.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2694 ( .DX(nn2694), .F0(nn2640), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_12|SUM_net ), .F3(dummy_abc_1679_) );
      defparam ii2694.CONFIG_DATA = 16'hB8B8;
      defparam ii2694.PLACE_LOCATION = "NONE";
      defparam ii2694.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2695 ( .DX(nn2695), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2694), .F2(dummy_abc_1680_), .F3(dummy_abc_1681_) );
      defparam ii2695.CONFIG_DATA = 16'h9999;
      defparam ii2695.PLACE_LOCATION = "NONE";
      defparam ii2695.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2696 ( .DX(nn2696), .F0(nn2641), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_13|SUM_net ), .F3(dummy_abc_1682_) );
      defparam ii2696.CONFIG_DATA = 16'hB8B8;
      defparam ii2696.PLACE_LOCATION = "NONE";
      defparam ii2696.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2697 ( .DX(nn2697), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2696), .F2(dummy_abc_1683_), .F3(dummy_abc_1684_) );
      defparam ii2697.CONFIG_DATA = 16'h9999;
      defparam ii2697.PLACE_LOCATION = "NONE";
      defparam ii2697.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2698 ( .DX(nn2698), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2678), .F2(dummy_abc_1685_), .F3(dummy_abc_1686_) );
      defparam ii2698.CONFIG_DATA = 16'h9999;
      defparam ii2698.PLACE_LOCATION = "NONE";
      defparam ii2698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2699 ( .DX(nn2699), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1687_), .F2(dummy_abc_1688_), .F3(dummy_abc_1689_) );
      defparam ii2699.CONFIG_DATA = 16'h5555;
      defparam ii2699.PLACE_LOCATION = "NONE";
      defparam ii2699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2700 ( .DX(nn2700), .F0(dummy_abc_1690_), .F1(dummy_abc_1691_), .F2(dummy_abc_1692_), .F3(dummy_abc_1693_) );
      defparam ii2700.CONFIG_DATA = 16'hFFFF;
      defparam ii2700.PLACE_LOCATION = "NONE";
      defparam ii2700.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_275_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_812_ ), 
        .DX( {nn2700, nn2699, nn2698, nn2697, nn2695, nn2693, nn2691, nn2689, 
              nn2688, nn2687, nn2686, nn2685, nn2684, nn2683, nn2682, nn2681, 
              nn2680, nn2679} ), 
        .SUM( {\coefcal1_divide_inst2_u148_XORCI_17|SUM_net , dummy_813_, 
              dummy_814_, dummy_815_, dummy_816_, dummy_817_, dummy_818_, dummy_819_, 
              dummy_820_, dummy_821_, dummy_822_, dummy_823_, dummy_824_, dummy_825_, 
              dummy_826_, dummy_827_, dummy_828_, dummy_829_} )
      );
    CS_LUT4_PRIM ii2721 ( .DX(nn2721), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_793_), .F3(dummy_abc_1694_) );
      defparam ii2721.CONFIG_DATA = 16'hA6A6;
      defparam ii2721.PLACE_LOCATION = "NONE";
      defparam ii2721.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2722 ( .DX(nn2722), .F0(dummy_793_), .F1(nn2629), .F2(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ), .F3(dummy_abc_1695_) );
      defparam ii2722.CONFIG_DATA = 16'hD8D8;
      defparam ii2722.PLACE_LOCATION = "NONE";
      defparam ii2722.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2723 ( .DX(nn2723), .F0(nn2630), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ), .F3(dummy_abc_1696_) );
      defparam ii2723.CONFIG_DATA = 16'hB8B8;
      defparam ii2723.PLACE_LOCATION = "NONE";
      defparam ii2723.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2724 ( .DX(nn2724), .F0(nn2631), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ), .F3(dummy_abc_1697_) );
      defparam ii2724.CONFIG_DATA = 16'hB8B8;
      defparam ii2724.PLACE_LOCATION = "NONE";
      defparam ii2724.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2725 ( .DX(nn2725), .F0(nn2632), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ), .F3(dummy_abc_1698_) );
      defparam ii2725.CONFIG_DATA = 16'hB8B8;
      defparam ii2725.PLACE_LOCATION = "NONE";
      defparam ii2725.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2726 ( .DX(nn2726), .F0(nn2633), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ), .F3(dummy_abc_1699_) );
      defparam ii2726.CONFIG_DATA = 16'hB8B8;
      defparam ii2726.PLACE_LOCATION = "NONE";
      defparam ii2726.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2727 ( .DX(nn2727), .F0(nn2634), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ), .F3(dummy_abc_1700_) );
      defparam ii2727.CONFIG_DATA = 16'hB8B8;
      defparam ii2727.PLACE_LOCATION = "NONE";
      defparam ii2727.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2728 ( .DX(nn2728), .F0(nn2635), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ), .F3(dummy_abc_1701_) );
      defparam ii2728.CONFIG_DATA = 16'hB8B8;
      defparam ii2728.PLACE_LOCATION = "NONE";
      defparam ii2728.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2729 ( .DX(nn2729), .F0(nn2636), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ), .F3(dummy_abc_1702_) );
      defparam ii2729.CONFIG_DATA = 16'hB8B8;
      defparam ii2729.PLACE_LOCATION = "NONE";
      defparam ii2729.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2730 ( .DX(nn2730), .F0(nn2637), .F1(dummy_793_), .F2(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ), .F3(dummy_abc_1703_) );
      defparam ii2730.CONFIG_DATA = 16'hB8B8;
      defparam ii2730.PLACE_LOCATION = "NONE";
      defparam ii2730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2731 ( .DX(nn2731), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1704_), .F3(dummy_abc_1705_) );
      defparam ii2731.CONFIG_DATA = 16'h9999;
      defparam ii2731.PLACE_LOCATION = "NONE";
      defparam ii2731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2732 ( .DX(nn2732), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_793_) );
      defparam ii2732.CONFIG_DATA = 16'hA569;
      defparam ii2732.PLACE_LOCATION = "NONE";
      defparam ii2732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2733 ( .DX(nn2733), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_793_), .F2(nn2629), .F3(\coefcal1_divide_inst2_u115_XORCI_1|SUM_net ) );
      defparam ii2733.CONFIG_DATA = 16'hA695;
      defparam ii2733.PLACE_LOCATION = "NONE";
      defparam ii2733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2734 ( .DX(nn2734), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2630), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_2|SUM_net ) );
      defparam ii2734.CONFIG_DATA = 16'h9A95;
      defparam ii2734.PLACE_LOCATION = "NONE";
      defparam ii2734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2735 ( .DX(nn2735), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2631), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_3|SUM_net ) );
      defparam ii2735.CONFIG_DATA = 16'h9A95;
      defparam ii2735.PLACE_LOCATION = "NONE";
      defparam ii2735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2736 ( .DX(nn2736), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2632), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_4|SUM_net ) );
      defparam ii2736.CONFIG_DATA = 16'h9A95;
      defparam ii2736.PLACE_LOCATION = "NONE";
      defparam ii2736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2737 ( .DX(nn2737), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2633), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_5|SUM_net ) );
      defparam ii2737.CONFIG_DATA = 16'h9A95;
      defparam ii2737.PLACE_LOCATION = "NONE";
      defparam ii2737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2738 ( .DX(nn2738), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2634), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_6|SUM_net ) );
      defparam ii2738.CONFIG_DATA = 16'h9A95;
      defparam ii2738.PLACE_LOCATION = "NONE";
      defparam ii2738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2739 ( .DX(nn2739), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2635), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_7|SUM_net ) );
      defparam ii2739.CONFIG_DATA = 16'h9A95;
      defparam ii2739.PLACE_LOCATION = "NONE";
      defparam ii2739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2740 ( .DX(nn2740), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2636), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_8|SUM_net ) );
      defparam ii2740.CONFIG_DATA = 16'h9A95;
      defparam ii2740.PLACE_LOCATION = "NONE";
      defparam ii2740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2741 ( .DX(nn2741), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2637), .F2(dummy_793_), .F3(\coefcal1_divide_inst2_u115_XORCI_9|SUM_net ) );
      defparam ii2741.CONFIG_DATA = 16'h9A95;
      defparam ii2741.PLACE_LOCATION = "NONE";
      defparam ii2741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2742 ( .DX(nn2742), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2690), .F2(dummy_abc_1706_), .F3(dummy_abc_1707_) );
      defparam ii2742.CONFIG_DATA = 16'h9999;
      defparam ii2742.PLACE_LOCATION = "NONE";
      defparam ii2742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2743 ( .DX(nn2743), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2692), .F2(dummy_abc_1708_), .F3(dummy_abc_1709_) );
      defparam ii2743.CONFIG_DATA = 16'h9999;
      defparam ii2743.PLACE_LOCATION = "NONE";
      defparam ii2743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2744 ( .DX(nn2744), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2694), .F2(dummy_abc_1710_), .F3(dummy_abc_1711_) );
      defparam ii2744.CONFIG_DATA = 16'h9999;
      defparam ii2744.PLACE_LOCATION = "NONE";
      defparam ii2744.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2745 ( .DX(nn2745), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2696), .F2(dummy_abc_1712_), .F3(dummy_abc_1713_) );
      defparam ii2745.CONFIG_DATA = 16'h9999;
      defparam ii2745.PLACE_LOCATION = "NONE";
      defparam ii2745.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2746 ( .DX(nn2746), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2678), .F2(dummy_abc_1714_), .F3(dummy_abc_1715_) );
      defparam ii2746.CONFIG_DATA = 16'h9999;
      defparam ii2746.PLACE_LOCATION = "NONE";
      defparam ii2746.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2747 ( .DX(nn2747), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(dummy_abc_1716_), .F2(dummy_abc_1717_), .F3(dummy_abc_1718_) );
      defparam ii2747.CONFIG_DATA = 16'h5555;
      defparam ii2747.PLACE_LOCATION = "NONE";
      defparam ii2747.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_259_ ( 
        .CA( {a_acc_en_cal1_u137_mac, nn2678, nn2696, nn2694, nn2692, nn2690, 
              nn2730, nn2729, nn2728, nn2727, nn2726, nn2725, nn2724, nn2723, 
              nn2722, nn2721, \coefcal1_yDividend__reg[1]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_199_ ), 
        .DX( {nn2747, nn2746, nn2745, nn2744, nn2743, nn2742, nn2741, nn2740, 
              nn2739, nn2738, nn2737, nn2736, nn2735, nn2734, nn2733, nn2732, 
              nn2731} ), 
        .SUM( {dummy_200_, \coefcal1_divide_inst2_u116_XORCI_15|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_14|SUM_net , \coefcal1_divide_inst2_u116_XORCI_13|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_12|SUM_net , \coefcal1_divide_inst2_u116_XORCI_11|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_10|SUM_net , \coefcal1_divide_inst2_u116_XORCI_9|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_8|SUM_net , \coefcal1_divide_inst2_u116_XORCI_7|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_6|SUM_net , \coefcal1_divide_inst2_u116_XORCI_5|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_4|SUM_net , \coefcal1_divide_inst2_u116_XORCI_3|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_2|SUM_net , \coefcal1_divide_inst2_u116_XORCI_1|SUM_net , 
              \coefcal1_divide_inst2_u116_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2767 ( .DX(nn2767), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(nn2678), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_15|SUM_net ) );
      defparam ii2767.CONFIG_DATA = 16'h202A;
      defparam ii2767.PLACE_LOCATION = "NONE";
      defparam ii2767.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2768 ( .DX(nn2768), .F0(\coefcal1_yDividend__reg[16]|Q_net ), .F1(\coefcal1_yDivisor__reg[16]|Q_net ), .F2(nn2767), .F3(dummy_abc_1719_) );
      defparam ii2768.CONFIG_DATA = 16'h0D0D;
      defparam ii2768.PLACE_LOCATION = "NONE";
      defparam ii2768.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2769 ( .DX(nn2769), .F0(dummy_abc_1720_), .F1(dummy_abc_1721_), .F2(dummy_abc_1722_), .F3(dummy_abc_1723_) );
      defparam ii2769.CONFIG_DATA = 16'hFFFF;
      defparam ii2769.PLACE_LOCATION = "NONE";
      defparam ii2769.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_260_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDividend__reg[16]|Q_net , 
              \coefcal1_yDividend__reg[15]|Q_net , \coefcal1_yDividend__reg[14]|Q_net , 
              \coefcal1_yDividend__reg[13]|Q_net , \coefcal1_yDividend__reg[12]|Q_net , 
              \coefcal1_yDividend__reg[11]|Q_net , \coefcal1_yDividend__reg[10]|Q_net , 
              \coefcal1_yDividend__reg[9]|Q_net , \coefcal1_yDividend__reg[8]|Q_net , 
              \coefcal1_yDividend__reg[7]|Q_net , \coefcal1_yDividend__reg[6]|Q_net , 
              \coefcal1_yDividend__reg[5]|Q_net , \coefcal1_yDividend__reg[4]|Q_net , 
              \coefcal1_yDividend__reg[3]|Q_net , \coefcal1_yDividend__reg[2]|Q_net , 
              \coefcal1_yDividend__reg[1]|Q_net , \coefcal1_yDividend__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_527_ ), 
        .DX( {nn2769, nn2768, nn1536, nn1535, nn1534, nn1533, nn1532, nn1531, 
              nn1530, nn1529, nn1528, nn1527, nn1526, nn1525, nn1524, nn1523, 
              nn1522, nn1521} ), 
        .SUM( {\coefcal1_divide_inst2_u118_XORCI_17|SUM_net , dummy_528_, 
              dummy_529_, dummy_530_, dummy_531_, dummy_532_, dummy_533_, dummy_534_, 
              dummy_535_, dummy_536_, dummy_537_, dummy_538_, dummy_539_, dummy_540_, 
              dummy_541_, dummy_542_, dummy_543_, dummy_544_} )
      );
    CS_LUT4_PRIM ii2790 ( .DX(nn2790), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(\coefcal1_yDivisor__reg[15]|Q_net ), .F2(\coefcal1_yDivisor__reg[16]|Q_net ), .F3(\coefcal1_yDivisor__reg[1]|Q_net ) );
      defparam ii2790.CONFIG_DATA = 16'h0001;
      defparam ii2790.PLACE_LOCATION = "NONE";
      defparam ii2790.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2791 ( .DX(nn2791), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(\coefcal1_yDivisor__reg[11]|Q_net ), .F2(\coefcal1_yDivisor__reg[12]|Q_net ), .F3(nn2790) );
      defparam ii2791.CONFIG_DATA = 16'h0100;
      defparam ii2791.PLACE_LOCATION = "NONE";
      defparam ii2791.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2792 ( .DX(nn2792), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(\coefcal1_yDivisor__reg[7]|Q_net ), .F2(\coefcal1_yDivisor__reg[8]|Q_net ), .F3(\coefcal1_yDivisor__reg[9]|Q_net ) );
      defparam ii2792.CONFIG_DATA = 16'h0001;
      defparam ii2792.PLACE_LOCATION = "NONE";
      defparam ii2792.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2793 ( .DX(nn2793), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(\coefcal1_yDivisor__reg[2]|Q_net ), .F2(\coefcal1_yDivisor__reg[5]|Q_net ), .F3(nn2792) );
      defparam ii2793.CONFIG_DATA = 16'h0100;
      defparam ii2793.PLACE_LOCATION = "NONE";
      defparam ii2793.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2794 ( .DX(nn2794), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(\coefcal1_yDivisor__reg[4]|Q_net ), .F2(nn2791), .F3(nn2793) );
      defparam ii2794.CONFIG_DATA = 16'h1000;
      defparam ii2794.PLACE_LOCATION = "NONE";
      defparam ii2794.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2795 ( .DX(nn2795), .F0(\coefcal1_yDivisor__reg[0]|Q_net ), .F1(nn2794), .F2(dummy_abc_1724_), .F3(dummy_abc_1725_) );
      defparam ii2795.CONFIG_DATA = 16'h4444;
      defparam ii2795.PLACE_LOCATION = "NONE";
      defparam ii2795.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2796 ( .DX(nn2796), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(dummy_abc_1726_), .F3(dummy_abc_1727_) );
      defparam ii2796.CONFIG_DATA = 16'h9999;
      defparam ii2796.PLACE_LOCATION = "NONE";
      defparam ii2796.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2797 ( .DX(nn2797), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(\coefcal1_yDivisor__reg[0]|Q_net ), .F2(\coefcal1_yDivisor__reg[1]|Q_net ), .F3(dummy_812_) );
      defparam ii2797.CONFIG_DATA = 16'hA569;
      defparam ii2797.PLACE_LOCATION = "NONE";
      defparam ii2797.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2798 ( .DX(nn2798), .F0(\coefcal1_yDivisor__reg[2]|Q_net ), .F1(dummy_812_), .F2(nn2721), .F3(\coefcal1_divide_inst2_u116_XORCI_1|SUM_net ) );
      defparam ii2798.CONFIG_DATA = 16'hA695;
      defparam ii2798.PLACE_LOCATION = "NONE";
      defparam ii2798.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2799 ( .DX(nn2799), .F0(\coefcal1_yDivisor__reg[3]|Q_net ), .F1(nn2722), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_2|SUM_net ) );
      defparam ii2799.CONFIG_DATA = 16'h9A95;
      defparam ii2799.PLACE_LOCATION = "NONE";
      defparam ii2799.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2800 ( .DX(nn2800), .F0(\coefcal1_yDivisor__reg[4]|Q_net ), .F1(nn2723), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_3|SUM_net ) );
      defparam ii2800.CONFIG_DATA = 16'h9A95;
      defparam ii2800.PLACE_LOCATION = "NONE";
      defparam ii2800.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2801 ( .DX(nn2801), .F0(\coefcal1_yDivisor__reg[5]|Q_net ), .F1(nn2724), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_4|SUM_net ) );
      defparam ii2801.CONFIG_DATA = 16'h9A95;
      defparam ii2801.PLACE_LOCATION = "NONE";
      defparam ii2801.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2802 ( .DX(nn2802), .F0(\coefcal1_yDivisor__reg[6]|Q_net ), .F1(nn2725), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_5|SUM_net ) );
      defparam ii2802.CONFIG_DATA = 16'h9A95;
      defparam ii2802.PLACE_LOCATION = "NONE";
      defparam ii2802.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2803 ( .DX(nn2803), .F0(\coefcal1_yDivisor__reg[7]|Q_net ), .F1(nn2726), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_6|SUM_net ) );
      defparam ii2803.CONFIG_DATA = 16'h9A95;
      defparam ii2803.PLACE_LOCATION = "NONE";
      defparam ii2803.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2804 ( .DX(nn2804), .F0(\coefcal1_yDivisor__reg[8]|Q_net ), .F1(nn2727), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_7|SUM_net ) );
      defparam ii2804.CONFIG_DATA = 16'h9A95;
      defparam ii2804.PLACE_LOCATION = "NONE";
      defparam ii2804.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2805 ( .DX(nn2805), .F0(\coefcal1_yDivisor__reg[9]|Q_net ), .F1(nn2728), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_8|SUM_net ) );
      defparam ii2805.CONFIG_DATA = 16'h9A95;
      defparam ii2805.PLACE_LOCATION = "NONE";
      defparam ii2805.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2806 ( .DX(nn2806), .F0(\coefcal1_yDivisor__reg[10]|Q_net ), .F1(nn2729), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_9|SUM_net ) );
      defparam ii2806.CONFIG_DATA = 16'h9A95;
      defparam ii2806.PLACE_LOCATION = "NONE";
      defparam ii2806.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2807 ( .DX(nn2807), .F0(\coefcal1_yDivisor__reg[11]|Q_net ), .F1(nn2730), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_10|SUM_net ) );
      defparam ii2807.CONFIG_DATA = 16'h9A95;
      defparam ii2807.PLACE_LOCATION = "NONE";
      defparam ii2807.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2808 ( .DX(nn2808), .F0(\coefcal1_yDivisor__reg[12]|Q_net ), .F1(nn2690), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_11|SUM_net ) );
      defparam ii2808.CONFIG_DATA = 16'h9A95;
      defparam ii2808.PLACE_LOCATION = "NONE";
      defparam ii2808.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2809 ( .DX(nn2809), .F0(\coefcal1_yDivisor__reg[13]|Q_net ), .F1(nn2692), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_12|SUM_net ) );
      defparam ii2809.CONFIG_DATA = 16'h9A95;
      defparam ii2809.PLACE_LOCATION = "NONE";
      defparam ii2809.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2810 ( .DX(nn2810), .F0(\coefcal1_yDivisor__reg[14]|Q_net ), .F1(nn2694), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_13|SUM_net ) );
      defparam ii2810.CONFIG_DATA = 16'h9A95;
      defparam ii2810.PLACE_LOCATION = "NONE";
      defparam ii2810.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2811 ( .DX(nn2811), .F0(\coefcal1_yDivisor__reg[15]|Q_net ), .F1(nn2696), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_14|SUM_net ) );
      defparam ii2811.CONFIG_DATA = 16'h9A95;
      defparam ii2811.PLACE_LOCATION = "NONE";
      defparam ii2811.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2812 ( .DX(nn2812), .F0(\coefcal1_yDivisor__reg[16]|Q_net ), .F1(nn2678), .F2(dummy_812_), .F3(\coefcal1_divide_inst2_u116_XORCI_15|SUM_net ) );
      defparam ii2812.CONFIG_DATA = 16'h9A95;
      defparam ii2812.PLACE_LOCATION = "NONE";
      defparam ii2812.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2813 ( .DX(nn2813), .F0(dummy_abc_1728_), .F1(dummy_abc_1729_), .F2(dummy_abc_1730_), .F3(dummy_abc_1731_) );
      defparam ii2813.CONFIG_DATA = 16'hFFFF;
      defparam ii2813.PLACE_LOCATION = "NONE";
      defparam ii2813.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_276_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_yDivisor__reg[16]|Q_net , 
              \coefcal1_yDivisor__reg[15]|Q_net , \coefcal1_yDivisor__reg[14]|Q_net , 
              \coefcal1_yDivisor__reg[13]|Q_net , \coefcal1_yDivisor__reg[12]|Q_net , 
              \coefcal1_yDivisor__reg[11]|Q_net , \coefcal1_yDivisor__reg[10]|Q_net , 
              \coefcal1_yDivisor__reg[9]|Q_net , \coefcal1_yDivisor__reg[8]|Q_net , 
              \coefcal1_yDivisor__reg[7]|Q_net , \coefcal1_yDivisor__reg[6]|Q_net , 
              \coefcal1_yDivisor__reg[5]|Q_net , \coefcal1_yDivisor__reg[4]|Q_net , 
              \coefcal1_yDivisor__reg[3]|Q_net , \coefcal1_yDivisor__reg[2]|Q_net , 
              \coefcal1_yDivisor__reg[1]|Q_net , \coefcal1_yDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_831_ ), 
        .DX( {nn2813, nn2812, nn2811, nn2810, nn2809, nn2808, nn2807, nn2806, 
              nn2805, nn2804, nn2803, nn2802, nn2801, nn2800, nn2799, nn2798, 
              nn2797, nn2796} ), 
        .SUM( {\coefcal1_divide_inst2_u150_XORCI_17|SUM_net , dummy_832_, 
              dummy_833_, dummy_834_, dummy_835_, dummy_836_, dummy_837_, dummy_838_, 
              dummy_839_, dummy_840_, dummy_841_, dummy_842_, dummy_843_, dummy_844_, 
              dummy_845_, dummy_846_, dummy_847_, dummy_848_} )
      );
    CS_LUT4_PRIM ii2834 ( .DX(nn2834), .F0(\coefcal1_yDividend__reg[0]|Q_net ), .F1(dummy_831_), .F2(nn2794), .F3(dummy_abc_1732_) );
      defparam ii2834.CONFIG_DATA = 16'h5C5C;
      defparam ii2834.PLACE_LOCATION = "NONE";
      defparam ii2834.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2835 ( .DX(nn2835), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2834) );
      defparam ii2835.CONFIG_DATA = 16'hFFFB;
      defparam ii2835.PLACE_LOCATION = "NONE";
      defparam ii2835.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2836 ( .DX(nn2836), .F0(\cal1_v__reg[0]|Q_net ), .F1(nn2835), .F2(dummy_abc_1733_), .F3(dummy_abc_1734_) );
      defparam ii2836.CONFIG_DATA = 16'h6666;
      defparam ii2836.PLACE_LOCATION = "NONE";
      defparam ii2836.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2837 ( .DX(nn2837), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2834) );
      defparam ii2837.CONFIG_DATA = 16'hFFFB;
      defparam ii2837.PLACE_LOCATION = "NONE";
      defparam ii2837.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2838 ( .DX(nn2838), .F0(\coefcal1_yDividend__reg[1]|Q_net ), .F1(dummy_812_), .F2(nn2794), .F3(dummy_abc_1735_) );
      defparam ii2838.CONFIG_DATA = 16'h5C5C;
      defparam ii2838.PLACE_LOCATION = "NONE";
      defparam ii2838.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2839 ( .DX(nn2839), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2838) );
      defparam ii2839.CONFIG_DATA = 16'h0004;
      defparam ii2839.PLACE_LOCATION = "NONE";
      defparam ii2839.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2840 ( .DX(nn2840), .F0(\coefcal1_yDividend__reg[2]|Q_net ), .F1(dummy_793_), .F2(nn2794), .F3(dummy_abc_1736_) );
      defparam ii2840.CONFIG_DATA = 16'h5C5C;
      defparam ii2840.PLACE_LOCATION = "NONE";
      defparam ii2840.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2841 ( .DX(nn2841), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2840) );
      defparam ii2841.CONFIG_DATA = 16'h0004;
      defparam ii2841.PLACE_LOCATION = "NONE";
      defparam ii2841.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2842 ( .DX(nn2842), .F0(\coefcal1_yDividend__reg[3]|Q_net ), .F1(dummy_774_), .F2(nn2794), .F3(dummy_abc_1737_) );
      defparam ii2842.CONFIG_DATA = 16'h5C5C;
      defparam ii2842.PLACE_LOCATION = "NONE";
      defparam ii2842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2843 ( .DX(nn2843), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2842) );
      defparam ii2843.CONFIG_DATA = 16'h0004;
      defparam ii2843.PLACE_LOCATION = "NONE";
      defparam ii2843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2844 ( .DX(nn2844), .F0(\coefcal1_yDividend__reg[4]|Q_net ), .F1(dummy_755_), .F2(nn2794), .F3(dummy_abc_1738_) );
      defparam ii2844.CONFIG_DATA = 16'h5C5C;
      defparam ii2844.PLACE_LOCATION = "NONE";
      defparam ii2844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2845 ( .DX(nn2845), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2844) );
      defparam ii2845.CONFIG_DATA = 16'h0004;
      defparam ii2845.PLACE_LOCATION = "NONE";
      defparam ii2845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2846 ( .DX(nn2846), .F0(\coefcal1_yDividend__reg[5]|Q_net ), .F1(dummy_736_), .F2(nn2794), .F3(dummy_abc_1739_) );
      defparam ii2846.CONFIG_DATA = 16'h5C5C;
      defparam ii2846.PLACE_LOCATION = "NONE";
      defparam ii2846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2847 ( .DX(nn2847), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2846) );
      defparam ii2847.CONFIG_DATA = 16'h0004;
      defparam ii2847.PLACE_LOCATION = "NONE";
      defparam ii2847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2848 ( .DX(nn2848), .F0(\coefcal1_yDividend__reg[6]|Q_net ), .F1(dummy_717_), .F2(nn2794), .F3(dummy_abc_1740_) );
      defparam ii2848.CONFIG_DATA = 16'h5C5C;
      defparam ii2848.PLACE_LOCATION = "NONE";
      defparam ii2848.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2849 ( .DX(nn2849), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2848) );
      defparam ii2849.CONFIG_DATA = 16'h0004;
      defparam ii2849.PLACE_LOCATION = "NONE";
      defparam ii2849.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2850 ( .DX(nn2850), .F0(\coefcal1_yDividend__reg[7]|Q_net ), .F1(dummy_698_), .F2(nn2794), .F3(dummy_abc_1741_) );
      defparam ii2850.CONFIG_DATA = 16'h5C5C;
      defparam ii2850.PLACE_LOCATION = "NONE";
      defparam ii2850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2851 ( .DX(nn2851), .F0(rst), .F1(dummy_527_), .F2(nn2795), .F3(nn2850) );
      defparam ii2851.CONFIG_DATA = 16'h0004;
      defparam ii2851.PLACE_LOCATION = "NONE";
      defparam ii2851.PCK_LOCATION = "NONE";
    scaler_ipc_adder_8 carry_8_279_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_dinxy_cen_cal1_u137_mac} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_888_ ), 
        .DX( {nn2851, nn2849, nn2847, nn2845, nn2843, nn2841, nn2839, nn2837} ), 
        .SUM( {\coefcal1_u62_XORCI_7|SUM_net , \coefcal1_u62_XORCI_6|SUM_net , 
              \coefcal1_u62_XORCI_5|SUM_net , \coefcal1_u62_XORCI_4|SUM_net , 
              \coefcal1_u62_XORCI_3|SUM_net , \coefcal1_u62_XORCI_2|SUM_net , 
              \coefcal1_u62_XORCI_1|SUM_net , \coefcal1_u62_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2862 ( .DX(nn2862), .F0(\cal1_v__reg[1]|Q_net ), .F1(\coefcal1_u62_XORCI_1|SUM_net ), .F2(dummy_abc_1742_), .F3(dummy_abc_1743_) );
      defparam ii2862.CONFIG_DATA = 16'h6666;
      defparam ii2862.PLACE_LOCATION = "NONE";
      defparam ii2862.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2863 ( .DX(nn2863), .F0(\cal1_v__reg[2]|Q_net ), .F1(\coefcal1_u62_XORCI_2|SUM_net ), .F2(dummy_abc_1744_), .F3(dummy_abc_1745_) );
      defparam ii2863.CONFIG_DATA = 16'h6666;
      defparam ii2863.PLACE_LOCATION = "NONE";
      defparam ii2863.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2864 ( .DX(nn2864), .F0(\cal1_v__reg[3]|Q_net ), .F1(\coefcal1_u62_XORCI_3|SUM_net ), .F2(dummy_abc_1746_), .F3(dummy_abc_1747_) );
      defparam ii2864.CONFIG_DATA = 16'h6666;
      defparam ii2864.PLACE_LOCATION = "NONE";
      defparam ii2864.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2865 ( .DX(nn2865), .F0(\cal1_v__reg[4]|Q_net ), .F1(\coefcal1_u62_XORCI_4|SUM_net ), .F2(dummy_abc_1748_), .F3(dummy_abc_1749_) );
      defparam ii2865.CONFIG_DATA = 16'h6666;
      defparam ii2865.PLACE_LOCATION = "NONE";
      defparam ii2865.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2866 ( .DX(nn2866), .F0(\cal1_v__reg[5]|Q_net ), .F1(\coefcal1_u62_XORCI_5|SUM_net ), .F2(dummy_abc_1750_), .F3(dummy_abc_1751_) );
      defparam ii2866.CONFIG_DATA = 16'h6666;
      defparam ii2866.PLACE_LOCATION = "NONE";
      defparam ii2866.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2867 ( .DX(nn2867), .F0(\cal1_v__reg[6]|Q_net ), .F1(\coefcal1_u62_XORCI_6|SUM_net ), .F2(dummy_abc_1752_), .F3(dummy_abc_1753_) );
      defparam ii2867.CONFIG_DATA = 16'h6666;
      defparam ii2867.PLACE_LOCATION = "NONE";
      defparam ii2867.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2868 ( .DX(nn2868), .F0(\cal1_v__reg[7]|Q_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_abc_1754_), .F3(dummy_abc_1755_) );
      defparam ii2868.CONFIG_DATA = 16'h6666;
      defparam ii2868.PLACE_LOCATION = "NONE";
      defparam ii2868.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2869 ( .DX(nn2869), .F0(\cal1_v__reg[8]|Q_net ), .F1(dummy_abc_1756_), .F2(dummy_abc_1757_), .F3(dummy_abc_1758_) );
      defparam ii2869.CONFIG_DATA = 16'hAAAA;
      defparam ii2869.PLACE_LOCATION = "NONE";
      defparam ii2869.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2870 ( .DX(nn2870), .F0(\cal1_v__reg[9]|Q_net ), .F1(dummy_abc_1759_), .F2(dummy_abc_1760_), .F3(dummy_abc_1761_) );
      defparam ii2870.CONFIG_DATA = 16'hAAAA;
      defparam ii2870.PLACE_LOCATION = "NONE";
      defparam ii2870.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2871 ( .DX(nn2871), .F0(\cal1_v__reg[10]|Q_net ), .F1(dummy_abc_1762_), .F2(dummy_abc_1763_), .F3(dummy_abc_1764_) );
      defparam ii2871.CONFIG_DATA = 16'hAAAA;
      defparam ii2871.PLACE_LOCATION = "NONE";
      defparam ii2871.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2872 ( .DX(nn2872), .F0(\cal1_v__reg[11]|Q_net ), .F1(dummy_abc_1765_), .F2(dummy_abc_1766_), .F3(dummy_abc_1767_) );
      defparam ii2872.CONFIG_DATA = 16'hAAAA;
      defparam ii2872.PLACE_LOCATION = "NONE";
      defparam ii2872.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2873 ( .DX(nn2873), .F0(\cal1_v__reg[12]|Q_net ), .F1(dummy_abc_1768_), .F2(dummy_abc_1769_), .F3(dummy_abc_1770_) );
      defparam ii2873.CONFIG_DATA = 16'hAAAA;
      defparam ii2873.PLACE_LOCATION = "NONE";
      defparam ii2873.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2874 ( .DX(nn2874), .F0(\cal1_v__reg[13]|Q_net ), .F1(dummy_abc_1771_), .F2(dummy_abc_1772_), .F3(dummy_abc_1773_) );
      defparam ii2874.CONFIG_DATA = 16'hAAAA;
      defparam ii2874.PLACE_LOCATION = "NONE";
      defparam ii2874.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2875 ( .DX(nn2875), .F0(\cal1_v__reg[14]|Q_net ), .F1(dummy_abc_1774_), .F2(dummy_abc_1775_), .F3(dummy_abc_1776_) );
      defparam ii2875.CONFIG_DATA = 16'hAAAA;
      defparam ii2875.PLACE_LOCATION = "NONE";
      defparam ii2875.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2876 ( .DX(nn2876), .F0(\cal1_v__reg[15]|Q_net ), .F1(dummy_abc_1777_), .F2(dummy_abc_1778_), .F3(dummy_abc_1779_) );
      defparam ii2876.CONFIG_DATA = 16'hAAAA;
      defparam ii2876.PLACE_LOCATION = "NONE";
      defparam ii2876.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2877 ( .DX(nn2877), .F0(\cal1_v__reg[16]|Q_net ), .F1(dummy_abc_1780_), .F2(dummy_abc_1781_), .F3(dummy_abc_1782_) );
      defparam ii2877.CONFIG_DATA = 16'hAAAA;
      defparam ii2877.PLACE_LOCATION = "NONE";
      defparam ii2877.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_198_ ( 
        .CA( {\cal1_v__reg[16]|Q_net , \cal1_v__reg[15]|Q_net , 
              \cal1_v__reg[14]|Q_net , \cal1_v__reg[13]|Q_net , \cal1_v__reg[12]|Q_net , 
              \cal1_v__reg[11]|Q_net , \cal1_v__reg[10]|Q_net , \cal1_v__reg[9]|Q_net , 
              \cal1_v__reg[8]|Q_net , \cal1_v__reg[7]|Q_net , \cal1_v__reg[6]|Q_net , 
              \cal1_v__reg[5]|Q_net , \cal1_v__reg[4]|Q_net , \cal1_v__reg[3]|Q_net , 
              \cal1_v__reg[2]|Q_net , \cal1_v__reg[1]|Q_net , \cal1_v__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_140_ ), 
        .DX( {nn2877, nn2876, nn2875, nn2874, nn2873, nn2872, nn2871, nn2870, 
              nn2869, nn2868, nn2867, nn2866, nn2865, nn2864, nn2863, nn2862, 
              nn2836} ), 
        .SUM( {\cal1_u128_XORCI_16|SUM_net , \cal1_u128_XORCI_15|SUM_net , 
              \cal1_u128_XORCI_14|SUM_net , \cal1_u128_XORCI_13|SUM_net , \cal1_u128_XORCI_12|SUM_net , 
              \cal1_u128_XORCI_11|SUM_net , \cal1_u128_XORCI_10|SUM_net , \cal1_u128_XORCI_9|SUM_net , 
              \cal1_u128_XORCI_8|SUM_net , \cal1_u128_XORCI_7|SUM_net , \cal1_u128_XORCI_6|SUM_net , 
              \cal1_u128_XORCI_5|SUM_net , \cal1_u128_XORCI_4|SUM_net , \cal1_u128_XORCI_3|SUM_net , 
              \cal1_u128_XORCI_2|SUM_net , \cal1_u128_XORCI_1|SUM_net , \cal1_u128_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2897 ( .DX(nn2897), .F0(\cal1_v__reg[6]|Q_net ), .F1(\cal1_v__reg[7]|Q_net ), .F2(\cal1_u128_XORCI_6|SUM_net ), .F3(\cal1_u128_XORCI_7|SUM_net ) );
      defparam ii2897.CONFIG_DATA = 16'h39C6;
      defparam ii2897.PLACE_LOCATION = "NONE";
      defparam ii2897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2898 ( .DX(nn2898), .F0(\cal1_v__reg[6]|Q_net ), .F1(\cal1_v__reg[7]|Q_net ), .F2(\cal1_u128_XORCI_6|SUM_net ), .F3(\cal1_u128_XORCI_7|SUM_net ) );
      defparam ii2898.CONFIG_DATA = 16'h08CE;
      defparam ii2898.PLACE_LOCATION = "NONE";
      defparam ii2898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2899 ( .DX(nn2899), .F0(\cal1_v__reg[8]|Q_net ), .F1(\cal1_u128_XORCI_8|SUM_net ), .F2(nn2897), .F3(nn2898) );
      defparam ii2899.CONFIG_DATA = 16'h0609;
      defparam ii2899.PLACE_LOCATION = "NONE";
      defparam ii2899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2900 ( .DX(nn2900), .F0(\cal1_v__reg[6]|Q_net ), .F1(dummy_62_), .F2(\cal1_u128_XORCI_6|SUM_net ), .F3(nn1517) );
      defparam ii2900.CONFIG_DATA = 16'h1200;
      defparam ii2900.PLACE_LOCATION = "NONE";
      defparam ii2900.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2901 ( .DX(nn2901), .F0(dummy_36_), .F1(nn1520), .F2(nn2899), .F3(nn2900) );
      defparam ii2901.CONFIG_DATA = 16'hF111;
      defparam ii2901.PLACE_LOCATION = "NONE";
      defparam ii2901.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2902 ( .DX(nn2902), .F0(dummy_62_), .F1(dummy_36_), .F2(dummy_23_), .F3(nn2899) );
      defparam ii2902.CONFIG_DATA = 16'h0004;
      defparam ii2902.PLACE_LOCATION = "NONE";
      defparam ii2902.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2903 ( .DX(nn2903), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1783_), .F3(dummy_abc_1784_) );
      defparam ii2903.CONFIG_DATA = 16'h9999;
      defparam ii2903.PLACE_LOCATION = "NONE";
      defparam ii2903.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2904 ( .DX(nn2904), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1785_), .F3(dummy_abc_1786_) );
      defparam ii2904.CONFIG_DATA = 16'h9999;
      defparam ii2904.PLACE_LOCATION = "NONE";
      defparam ii2904.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2905 ( .DX(nn2905), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_abc_1787_), .F3(dummy_abc_1788_) );
      defparam ii2905.CONFIG_DATA = 16'h9999;
      defparam ii2905.PLACE_LOCATION = "NONE";
      defparam ii2905.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2906 ( .DX(nn2906), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[3]|Q_net ), .F2(dummy_abc_1789_), .F3(dummy_abc_1790_) );
      defparam ii2906.CONFIG_DATA = 16'h9999;
      defparam ii2906.PLACE_LOCATION = "NONE";
      defparam ii2906.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2907 ( .DX(nn2907), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[4]|Q_net ), .F2(dummy_abc_1791_), .F3(dummy_abc_1792_) );
      defparam ii2907.CONFIG_DATA = 16'h9999;
      defparam ii2907.PLACE_LOCATION = "NONE";
      defparam ii2907.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2908 ( .DX(nn2908), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[5]|Q_net ), .F2(dummy_abc_1793_), .F3(dummy_abc_1794_) );
      defparam ii2908.CONFIG_DATA = 16'h9999;
      defparam ii2908.PLACE_LOCATION = "NONE";
      defparam ii2908.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2909 ( .DX(nn2909), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[6]|Q_net ), .F2(dummy_abc_1795_), .F3(dummy_abc_1796_) );
      defparam ii2909.CONFIG_DATA = 16'h9999;
      defparam ii2909.PLACE_LOCATION = "NONE";
      defparam ii2909.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2910 ( .DX(nn2910), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[7]|Q_net ), .F2(dummy_abc_1797_), .F3(dummy_abc_1798_) );
      defparam ii2910.CONFIG_DATA = 16'h9999;
      defparam ii2910.PLACE_LOCATION = "NONE";
      defparam ii2910.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2911 ( .DX(nn2911), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[8]|Q_net ), .F2(dummy_abc_1799_), .F3(dummy_abc_1800_) );
      defparam ii2911.CONFIG_DATA = 16'h9999;
      defparam ii2911.PLACE_LOCATION = "NONE";
      defparam ii2911.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2912 ( .DX(nn2912), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[9]|Q_net ), .F2(dummy_abc_1801_), .F3(dummy_abc_1802_) );
      defparam ii2912.CONFIG_DATA = 16'h9999;
      defparam ii2912.PLACE_LOCATION = "NONE";
      defparam ii2912.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2913 ( .DX(nn2913), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[10]|Q_net ), .F2(dummy_abc_1803_), .F3(dummy_abc_1804_) );
      defparam ii2913.CONFIG_DATA = 16'h9999;
      defparam ii2913.PLACE_LOCATION = "NONE";
      defparam ii2913.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2914 ( .DX(nn2914), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[11]|Q_net ), .F2(dummy_abc_1805_), .F3(dummy_abc_1806_) );
      defparam ii2914.CONFIG_DATA = 16'h9999;
      defparam ii2914.PLACE_LOCATION = "NONE";
      defparam ii2914.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2915 ( .DX(nn2915), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[12]|Q_net ), .F2(dummy_abc_1807_), .F3(dummy_abc_1808_) );
      defparam ii2915.CONFIG_DATA = 16'h9999;
      defparam ii2915.PLACE_LOCATION = "NONE";
      defparam ii2915.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2916 ( .DX(nn2916), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[13]|Q_net ), .F2(dummy_abc_1809_), .F3(dummy_abc_1810_) );
      defparam ii2916.CONFIG_DATA = 16'h9999;
      defparam ii2916.PLACE_LOCATION = "NONE";
      defparam ii2916.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2917 ( .DX(nn2917), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[14]|Q_net ), .F2(dummy_abc_1811_), .F3(dummy_abc_1812_) );
      defparam ii2917.CONFIG_DATA = 16'h9999;
      defparam ii2917.PLACE_LOCATION = "NONE";
      defparam ii2917.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2918 ( .DX(nn2918), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[15]|Q_net ), .F2(dummy_abc_1813_), .F3(dummy_abc_1814_) );
      defparam ii2918.CONFIG_DATA = 16'h9999;
      defparam ii2918.PLACE_LOCATION = "NONE";
      defparam ii2918.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2919 ( .DX(nn2919), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1815_), .F3(dummy_abc_1816_) );
      defparam ii2919.CONFIG_DATA = 16'h9999;
      defparam ii2919.PLACE_LOCATION = "NONE";
      defparam ii2919.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2920 ( .DX(nn2920), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1817_), .F3(dummy_abc_1818_) );
      defparam ii2920.CONFIG_DATA = 16'h9999;
      defparam ii2920.PLACE_LOCATION = "NONE";
      defparam ii2920.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2921 ( .DX(nn2921), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1819_), .F3(dummy_abc_1820_) );
      defparam ii2921.CONFIG_DATA = 16'h9999;
      defparam ii2921.PLACE_LOCATION = "NONE";
      defparam ii2921.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2922 ( .DX(nn2922), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_abc_1821_), .F2(dummy_abc_1822_), .F3(dummy_abc_1823_) );
      defparam ii2922.CONFIG_DATA = 16'h5555;
      defparam ii2922.PLACE_LOCATION = "NONE";
      defparam ii2922.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2923 ( .DX(nn2923), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1824_), .F2(dummy_abc_1825_), .F3(dummy_abc_1826_) );
      defparam ii2923.CONFIG_DATA = 16'h5555;
      defparam ii2923.PLACE_LOCATION = "NONE";
      defparam ii2923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2924 ( .DX(nn2924), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1827_), .F2(dummy_abc_1828_), .F3(dummy_abc_1829_) );
      defparam ii2924.CONFIG_DATA = 16'h5555;
      defparam ii2924.PLACE_LOCATION = "NONE";
      defparam ii2924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2925 ( .DX(nn2925), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1830_), .F2(dummy_abc_1831_), .F3(dummy_abc_1832_) );
      defparam ii2925.CONFIG_DATA = 16'h5555;
      defparam ii2925.PLACE_LOCATION = "NONE";
      defparam ii2925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2926 ( .DX(nn2926), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1833_), .F2(dummy_abc_1834_), .F3(dummy_abc_1835_) );
      defparam ii2926.CONFIG_DATA = 16'h5555;
      defparam ii2926.PLACE_LOCATION = "NONE";
      defparam ii2926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2927 ( .DX(nn2927), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1836_), .F2(dummy_abc_1837_), .F3(dummy_abc_1838_) );
      defparam ii2927.CONFIG_DATA = 16'h5555;
      defparam ii2927.PLACE_LOCATION = "NONE";
      defparam ii2927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2928 ( .DX(nn2928), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1839_), .F2(dummy_abc_1840_), .F3(dummy_abc_1841_) );
      defparam ii2928.CONFIG_DATA = 16'h5555;
      defparam ii2928.PLACE_LOCATION = "NONE";
      defparam ii2928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2929 ( .DX(nn2929), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1842_), .F2(dummy_abc_1843_), .F3(dummy_abc_1844_) );
      defparam ii2929.CONFIG_DATA = 16'h5555;
      defparam ii2929.PLACE_LOCATION = "NONE";
      defparam ii2929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2930 ( .DX(nn2930), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1845_), .F2(dummy_abc_1846_), .F3(dummy_abc_1847_) );
      defparam ii2930.CONFIG_DATA = 16'h5555;
      defparam ii2930.PLACE_LOCATION = "NONE";
      defparam ii2930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2931 ( .DX(nn2931), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1848_), .F2(dummy_abc_1849_), .F3(dummy_abc_1850_) );
      defparam ii2931.CONFIG_DATA = 16'h5555;
      defparam ii2931.PLACE_LOCATION = "NONE";
      defparam ii2931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2932 ( .DX(nn2932), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1851_), .F2(dummy_abc_1852_), .F3(dummy_abc_1853_) );
      defparam ii2932.CONFIG_DATA = 16'h5555;
      defparam ii2932.PLACE_LOCATION = "NONE";
      defparam ii2932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2933 ( .DX(nn2933), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1854_), .F2(dummy_abc_1855_), .F3(dummy_abc_1856_) );
      defparam ii2933.CONFIG_DATA = 16'h5555;
      defparam ii2933.PLACE_LOCATION = "NONE";
      defparam ii2933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2934 ( .DX(nn2934), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1857_), .F2(dummy_abc_1858_), .F3(dummy_abc_1859_) );
      defparam ii2934.CONFIG_DATA = 16'h5555;
      defparam ii2934.PLACE_LOCATION = "NONE";
      defparam ii2934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2935 ( .DX(nn2935), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1860_), .F2(dummy_abc_1861_), .F3(dummy_abc_1862_) );
      defparam ii2935.CONFIG_DATA = 16'h5555;
      defparam ii2935.PLACE_LOCATION = "NONE";
      defparam ii2935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2936 ( .DX(nn2936), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1863_), .F2(dummy_abc_1864_), .F3(dummy_abc_1865_) );
      defparam ii2936.CONFIG_DATA = 16'h5555;
      defparam ii2936.PLACE_LOCATION = "NONE";
      defparam ii2936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2937 ( .DX(nn2937), .F0(dummy_abc_1866_), .F1(dummy_abc_1867_), .F2(dummy_abc_1868_), .F3(dummy_abc_1869_) );
      defparam ii2937.CONFIG_DATA = 16'hFFFF;
      defparam ii2937.PLACE_LOCATION = "NONE";
      defparam ii2937.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_229_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_223_ ), 
        .DX( {nn2937, nn2936, nn2935, nn2934, nn2933, nn2932, nn2931, nn2930, 
              nn2929, nn2928, nn2927, nn2926, nn2925, nn2924, nn2923, nn2922, 
              nn2921, nn2920} ), 
        .SUM( {\coefcal1_divide_inst1_u120_XORCI_17|SUM_net , dummy_224_, 
              dummy_225_, dummy_226_, dummy_227_, dummy_228_, dummy_229_, dummy_230_, 
              dummy_231_, dummy_232_, dummy_233_, dummy_234_, dummy_235_, dummy_236_, 
              dummy_237_, dummy_238_, dummy_239_, dummy_240_} )
      );
    CS_LUT4_PRIM ii2958 ( .DX(nn2958), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_223_) );
      defparam ii2958.CONFIG_DATA = 16'hA569;
      defparam ii2958.PLACE_LOCATION = "NONE";
      defparam ii2958.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2959 ( .DX(nn2959), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1870_), .F3(dummy_abc_1871_) );
      defparam ii2959.CONFIG_DATA = 16'h9999;
      defparam ii2959.PLACE_LOCATION = "NONE";
      defparam ii2959.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2960 ( .DX(nn2960), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[1]|Q_net ), .F2(dummy_abc_1872_), .F3(dummy_abc_1873_) );
      defparam ii2960.CONFIG_DATA = 16'h9999;
      defparam ii2960.PLACE_LOCATION = "NONE";
      defparam ii2960.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2961 ( .DX(nn2961), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_abc_1874_), .F2(dummy_abc_1875_), .F3(dummy_abc_1876_) );
      defparam ii2961.CONFIG_DATA = 16'h5555;
      defparam ii2961.PLACE_LOCATION = "NONE";
      defparam ii2961.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2962 ( .DX(nn2962), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1877_), .F2(dummy_abc_1878_), .F3(dummy_abc_1879_) );
      defparam ii2962.CONFIG_DATA = 16'h5555;
      defparam ii2962.PLACE_LOCATION = "NONE";
      defparam ii2962.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2963 ( .DX(nn2963), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1880_), .F2(dummy_abc_1881_), .F3(dummy_abc_1882_) );
      defparam ii2963.CONFIG_DATA = 16'h5555;
      defparam ii2963.PLACE_LOCATION = "NONE";
      defparam ii2963.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2964 ( .DX(nn2964), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1883_), .F2(dummy_abc_1884_), .F3(dummy_abc_1885_) );
      defparam ii2964.CONFIG_DATA = 16'h5555;
      defparam ii2964.PLACE_LOCATION = "NONE";
      defparam ii2964.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2965 ( .DX(nn2965), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1886_), .F2(dummy_abc_1887_), .F3(dummy_abc_1888_) );
      defparam ii2965.CONFIG_DATA = 16'h5555;
      defparam ii2965.PLACE_LOCATION = "NONE";
      defparam ii2965.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2966 ( .DX(nn2966), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1889_), .F2(dummy_abc_1890_), .F3(dummy_abc_1891_) );
      defparam ii2966.CONFIG_DATA = 16'h5555;
      defparam ii2966.PLACE_LOCATION = "NONE";
      defparam ii2966.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2967 ( .DX(nn2967), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1892_), .F2(dummy_abc_1893_), .F3(dummy_abc_1894_) );
      defparam ii2967.CONFIG_DATA = 16'h5555;
      defparam ii2967.PLACE_LOCATION = "NONE";
      defparam ii2967.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2968 ( .DX(nn2968), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1895_), .F2(dummy_abc_1896_), .F3(dummy_abc_1897_) );
      defparam ii2968.CONFIG_DATA = 16'h5555;
      defparam ii2968.PLACE_LOCATION = "NONE";
      defparam ii2968.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2969 ( .DX(nn2969), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1898_), .F2(dummy_abc_1899_), .F3(dummy_abc_1900_) );
      defparam ii2969.CONFIG_DATA = 16'h5555;
      defparam ii2969.PLACE_LOCATION = "NONE";
      defparam ii2969.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2970 ( .DX(nn2970), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1901_), .F2(dummy_abc_1902_), .F3(dummy_abc_1903_) );
      defparam ii2970.CONFIG_DATA = 16'h5555;
      defparam ii2970.PLACE_LOCATION = "NONE";
      defparam ii2970.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2971 ( .DX(nn2971), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1904_), .F2(dummy_abc_1905_), .F3(dummy_abc_1906_) );
      defparam ii2971.CONFIG_DATA = 16'h5555;
      defparam ii2971.PLACE_LOCATION = "NONE";
      defparam ii2971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2972 ( .DX(nn2972), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1907_), .F2(dummy_abc_1908_), .F3(dummy_abc_1909_) );
      defparam ii2972.CONFIG_DATA = 16'h5555;
      defparam ii2972.PLACE_LOCATION = "NONE";
      defparam ii2972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2973 ( .DX(nn2973), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1910_), .F2(dummy_abc_1911_), .F3(dummy_abc_1912_) );
      defparam ii2973.CONFIG_DATA = 16'h5555;
      defparam ii2973.PLACE_LOCATION = "NONE";
      defparam ii2973.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2974 ( .DX(nn2974), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1913_), .F2(dummy_abc_1914_), .F3(dummy_abc_1915_) );
      defparam ii2974.CONFIG_DATA = 16'h5555;
      defparam ii2974.PLACE_LOCATION = "NONE";
      defparam ii2974.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2975 ( .DX(nn2975), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1916_), .F2(dummy_abc_1917_), .F3(dummy_abc_1918_) );
      defparam ii2975.CONFIG_DATA = 16'h5555;
      defparam ii2975.PLACE_LOCATION = "NONE";
      defparam ii2975.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_214_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, \coefcal1_xDividend__reg[16]|Q_net , 
              \coefcal1_xDividend__reg[15]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_141_ ), 
        .DX( {nn2975, nn2974, nn2973, nn2972, nn2971, nn2970, nn2969, nn2968, 
              nn2967, nn2966, nn2965, nn2964, nn2963, nn2962, nn2961, nn2960, 
              nn2959} ), 
        .SUM( {dummy_142_, \coefcal1_divide_inst1_u102_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_14|SUM_net , \coefcal1_divide_inst1_u102_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_12|SUM_net , \coefcal1_divide_inst1_u102_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_10|SUM_net , \coefcal1_divide_inst1_u102_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_8|SUM_net , \coefcal1_divide_inst1_u102_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_6|SUM_net , \coefcal1_divide_inst1_u102_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_4|SUM_net , \coefcal1_divide_inst1_u102_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_2|SUM_net , \coefcal1_divide_inst1_u102_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u102_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii2995 ( .DX(nn2995), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_223_), .F3(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ) );
      defparam ii2995.CONFIG_DATA = 16'h9C93;
      defparam ii2995.PLACE_LOCATION = "NONE";
      defparam ii2995.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2996 ( .DX(nn2996), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1919_), .F2(dummy_abc_1920_), .F3(dummy_abc_1921_) );
      defparam ii2996.CONFIG_DATA = 16'h5555;
      defparam ii2996.PLACE_LOCATION = "NONE";
      defparam ii2996.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2997 ( .DX(nn2997), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1922_), .F2(dummy_abc_1923_), .F3(dummy_abc_1924_) );
      defparam ii2997.CONFIG_DATA = 16'h5555;
      defparam ii2997.PLACE_LOCATION = "NONE";
      defparam ii2997.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2998 ( .DX(nn2998), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1925_), .F2(dummy_abc_1926_), .F3(dummy_abc_1927_) );
      defparam ii2998.CONFIG_DATA = 16'h5555;
      defparam ii2998.PLACE_LOCATION = "NONE";
      defparam ii2998.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii2999 ( .DX(nn2999), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1928_), .F2(dummy_abc_1929_), .F3(dummy_abc_1930_) );
      defparam ii2999.CONFIG_DATA = 16'h5555;
      defparam ii2999.PLACE_LOCATION = "NONE";
      defparam ii2999.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3000 ( .DX(nn3000), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1931_), .F2(dummy_abc_1932_), .F3(dummy_abc_1933_) );
      defparam ii3000.CONFIG_DATA = 16'h5555;
      defparam ii3000.PLACE_LOCATION = "NONE";
      defparam ii3000.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3001 ( .DX(nn3001), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1934_), .F2(dummy_abc_1935_), .F3(dummy_abc_1936_) );
      defparam ii3001.CONFIG_DATA = 16'h5555;
      defparam ii3001.PLACE_LOCATION = "NONE";
      defparam ii3001.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3002 ( .DX(nn3002), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1937_), .F2(dummy_abc_1938_), .F3(dummy_abc_1939_) );
      defparam ii3002.CONFIG_DATA = 16'h5555;
      defparam ii3002.PLACE_LOCATION = "NONE";
      defparam ii3002.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3003 ( .DX(nn3003), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1940_), .F2(dummy_abc_1941_), .F3(dummy_abc_1942_) );
      defparam ii3003.CONFIG_DATA = 16'h5555;
      defparam ii3003.PLACE_LOCATION = "NONE";
      defparam ii3003.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3004 ( .DX(nn3004), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1943_), .F2(dummy_abc_1944_), .F3(dummy_abc_1945_) );
      defparam ii3004.CONFIG_DATA = 16'h5555;
      defparam ii3004.PLACE_LOCATION = "NONE";
      defparam ii3004.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3005 ( .DX(nn3005), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1946_), .F2(dummy_abc_1947_), .F3(dummy_abc_1948_) );
      defparam ii3005.CONFIG_DATA = 16'h5555;
      defparam ii3005.PLACE_LOCATION = "NONE";
      defparam ii3005.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3006 ( .DX(nn3006), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_1949_), .F2(dummy_abc_1950_), .F3(dummy_abc_1951_) );
      defparam ii3006.CONFIG_DATA = 16'h5555;
      defparam ii3006.PLACE_LOCATION = "NONE";
      defparam ii3006.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3007 ( .DX(nn3007), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_1952_), .F2(dummy_abc_1953_), .F3(dummy_abc_1954_) );
      defparam ii3007.CONFIG_DATA = 16'h5555;
      defparam ii3007.PLACE_LOCATION = "NONE";
      defparam ii3007.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3008 ( .DX(nn3008), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_1955_), .F2(dummy_abc_1956_), .F3(dummy_abc_1957_) );
      defparam ii3008.CONFIG_DATA = 16'h5555;
      defparam ii3008.PLACE_LOCATION = "NONE";
      defparam ii3008.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3009 ( .DX(nn3009), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_1958_), .F2(dummy_abc_1959_), .F3(dummy_abc_1960_) );
      defparam ii3009.CONFIG_DATA = 16'h5555;
      defparam ii3009.PLACE_LOCATION = "NONE";
      defparam ii3009.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3010 ( .DX(nn3010), .F0(dummy_abc_1961_), .F1(dummy_abc_1962_), .F2(dummy_abc_1963_), .F3(dummy_abc_1964_) );
      defparam ii3010.CONFIG_DATA = 16'hFFFF;
      defparam ii3010.PLACE_LOCATION = "NONE";
      defparam ii3010.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_230_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_242_ ), 
        .DX( {nn3010, nn3009, nn3008, nn3007, nn3006, nn3005, nn3004, nn3003, 
              nn3002, nn3001, nn3000, nn2999, nn2998, nn2997, nn2996, nn2995, 
              nn2958, nn2919} ), 
        .SUM( {\coefcal1_divide_inst1_u122_XORCI_17|SUM_net , dummy_243_, 
              dummy_244_, dummy_245_, dummy_246_, dummy_247_, dummy_248_, dummy_249_, 
              dummy_250_, dummy_251_, dummy_252_, dummy_253_, dummy_254_, dummy_255_, 
              dummy_256_, dummy_257_, dummy_258_, dummy_259_} )
      );
    CS_LUT4_PRIM ii3031 ( .DX(nn3031), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1965_), .F3(dummy_abc_1966_) );
      defparam ii3031.CONFIG_DATA = 16'h9999;
      defparam ii3031.PLACE_LOCATION = "NONE";
      defparam ii3031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3032 ( .DX(nn3032), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_242_) );
      defparam ii3032.CONFIG_DATA = 16'hA569;
      defparam ii3032.PLACE_LOCATION = "NONE";
      defparam ii3032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3033 ( .DX(nn3033), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_223_), .F3(dummy_abc_1967_) );
      defparam ii3033.CONFIG_DATA = 16'hA6A6;
      defparam ii3033.PLACE_LOCATION = "NONE";
      defparam ii3033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3034 ( .DX(nn3034), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(dummy_223_), .F2(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ), .F3(dummy_abc_1968_) );
      defparam ii3034.CONFIG_DATA = 16'hB8B8;
      defparam ii3034.PLACE_LOCATION = "NONE";
      defparam ii3034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3035 ( .DX(nn3035), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_1969_), .F3(dummy_abc_1970_) );
      defparam ii3035.CONFIG_DATA = 16'h9999;
      defparam ii3035.PLACE_LOCATION = "NONE";
      defparam ii3035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3036 ( .DX(nn3036), .F0(\coefcal1_xDividend__reg[15]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_223_) );
      defparam ii3036.CONFIG_DATA = 16'hA569;
      defparam ii3036.PLACE_LOCATION = "NONE";
      defparam ii3036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3037 ( .DX(nn3037), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(dummy_223_), .F3(\coefcal1_divide_inst1_u102_XORCI_1|SUM_net ) );
      defparam ii3037.CONFIG_DATA = 16'h9C93;
      defparam ii3037.PLACE_LOCATION = "NONE";
      defparam ii3037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3038 ( .DX(nn3038), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(dummy_abc_1971_), .F2(dummy_abc_1972_), .F3(dummy_abc_1973_) );
      defparam ii3038.CONFIG_DATA = 16'h5555;
      defparam ii3038.PLACE_LOCATION = "NONE";
      defparam ii3038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3039 ( .DX(nn3039), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_1974_), .F2(dummy_abc_1975_), .F3(dummy_abc_1976_) );
      defparam ii3039.CONFIG_DATA = 16'h5555;
      defparam ii3039.PLACE_LOCATION = "NONE";
      defparam ii3039.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3040 ( .DX(nn3040), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_1977_), .F2(dummy_abc_1978_), .F3(dummy_abc_1979_) );
      defparam ii3040.CONFIG_DATA = 16'h5555;
      defparam ii3040.PLACE_LOCATION = "NONE";
      defparam ii3040.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3041 ( .DX(nn3041), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_1980_), .F2(dummy_abc_1981_), .F3(dummy_abc_1982_) );
      defparam ii3041.CONFIG_DATA = 16'h5555;
      defparam ii3041.PLACE_LOCATION = "NONE";
      defparam ii3041.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3042 ( .DX(nn3042), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_1983_), .F2(dummy_abc_1984_), .F3(dummy_abc_1985_) );
      defparam ii3042.CONFIG_DATA = 16'h5555;
      defparam ii3042.PLACE_LOCATION = "NONE";
      defparam ii3042.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3043 ( .DX(nn3043), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_1986_), .F2(dummy_abc_1987_), .F3(dummy_abc_1988_) );
      defparam ii3043.CONFIG_DATA = 16'h5555;
      defparam ii3043.PLACE_LOCATION = "NONE";
      defparam ii3043.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3044 ( .DX(nn3044), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_1989_), .F2(dummy_abc_1990_), .F3(dummy_abc_1991_) );
      defparam ii3044.CONFIG_DATA = 16'h5555;
      defparam ii3044.PLACE_LOCATION = "NONE";
      defparam ii3044.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3045 ( .DX(nn3045), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_1992_), .F2(dummy_abc_1993_), .F3(dummy_abc_1994_) );
      defparam ii3045.CONFIG_DATA = 16'h5555;
      defparam ii3045.PLACE_LOCATION = "NONE";
      defparam ii3045.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3046 ( .DX(nn3046), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_1995_), .F2(dummy_abc_1996_), .F3(dummy_abc_1997_) );
      defparam ii3046.CONFIG_DATA = 16'h5555;
      defparam ii3046.PLACE_LOCATION = "NONE";
      defparam ii3046.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3047 ( .DX(nn3047), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_1998_), .F2(dummy_abc_1999_), .F3(dummy_abc_2000_) );
      defparam ii3047.CONFIG_DATA = 16'h5555;
      defparam ii3047.PLACE_LOCATION = "NONE";
      defparam ii3047.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3048 ( .DX(nn3048), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2001_), .F2(dummy_abc_2002_), .F3(dummy_abc_2003_) );
      defparam ii3048.CONFIG_DATA = 16'h5555;
      defparam ii3048.PLACE_LOCATION = "NONE";
      defparam ii3048.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3049 ( .DX(nn3049), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2004_), .F2(dummy_abc_2005_), .F3(dummy_abc_2006_) );
      defparam ii3049.CONFIG_DATA = 16'h5555;
      defparam ii3049.PLACE_LOCATION = "NONE";
      defparam ii3049.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3050 ( .DX(nn3050), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2007_), .F2(dummy_abc_2008_), .F3(dummy_abc_2009_) );
      defparam ii3050.CONFIG_DATA = 16'h5555;
      defparam ii3050.PLACE_LOCATION = "NONE";
      defparam ii3050.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3051 ( .DX(nn3051), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2010_), .F2(dummy_abc_2011_), .F3(dummy_abc_2012_) );
      defparam ii3051.CONFIG_DATA = 16'h5555;
      defparam ii3051.PLACE_LOCATION = "NONE";
      defparam ii3051.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_215_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3034, 
              nn3033, \coefcal1_xDividend__reg[14]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_143_ ), 
        .DX( {nn3051, nn3050, nn3049, nn3048, nn3047, nn3046, nn3045, nn3044, 
              nn3043, nn3042, nn3041, nn3040, nn3039, nn3038, nn3037, nn3036, 
              nn3035} ), 
        .SUM( {dummy_144_, \coefcal1_divide_inst1_u103_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_14|SUM_net , \coefcal1_divide_inst1_u103_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_12|SUM_net , \coefcal1_divide_inst1_u103_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_10|SUM_net , \coefcal1_divide_inst1_u103_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_8|SUM_net , \coefcal1_divide_inst1_u103_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_6|SUM_net , \coefcal1_divide_inst1_u103_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_4|SUM_net , \coefcal1_divide_inst1_u103_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_2|SUM_net , \coefcal1_divide_inst1_u103_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u103_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3071 ( .DX(nn3071), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_242_), .F2(nn3033), .F3(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ) );
      defparam ii3071.CONFIG_DATA = 16'hA695;
      defparam ii3071.PLACE_LOCATION = "NONE";
      defparam ii3071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3072 ( .DX(nn3072), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3034), .F2(dummy_242_), .F3(\coefcal1_divide_inst1_u103_XORCI_2|SUM_net ) );
      defparam ii3072.CONFIG_DATA = 16'h9A95;
      defparam ii3072.PLACE_LOCATION = "NONE";
      defparam ii3072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3073 ( .DX(nn3073), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_2013_), .F2(dummy_abc_2014_), .F3(dummy_abc_2015_) );
      defparam ii3073.CONFIG_DATA = 16'h5555;
      defparam ii3073.PLACE_LOCATION = "NONE";
      defparam ii3073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3074 ( .DX(nn3074), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_2016_), .F2(dummy_abc_2017_), .F3(dummy_abc_2018_) );
      defparam ii3074.CONFIG_DATA = 16'h5555;
      defparam ii3074.PLACE_LOCATION = "NONE";
      defparam ii3074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3075 ( .DX(nn3075), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2019_), .F2(dummy_abc_2020_), .F3(dummy_abc_2021_) );
      defparam ii3075.CONFIG_DATA = 16'h5555;
      defparam ii3075.PLACE_LOCATION = "NONE";
      defparam ii3075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3076 ( .DX(nn3076), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2022_), .F2(dummy_abc_2023_), .F3(dummy_abc_2024_) );
      defparam ii3076.CONFIG_DATA = 16'h5555;
      defparam ii3076.PLACE_LOCATION = "NONE";
      defparam ii3076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3077 ( .DX(nn3077), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2025_), .F2(dummy_abc_2026_), .F3(dummy_abc_2027_) );
      defparam ii3077.CONFIG_DATA = 16'h5555;
      defparam ii3077.PLACE_LOCATION = "NONE";
      defparam ii3077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3078 ( .DX(nn3078), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2028_), .F2(dummy_abc_2029_), .F3(dummy_abc_2030_) );
      defparam ii3078.CONFIG_DATA = 16'h5555;
      defparam ii3078.PLACE_LOCATION = "NONE";
      defparam ii3078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3079 ( .DX(nn3079), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2031_), .F2(dummy_abc_2032_), .F3(dummy_abc_2033_) );
      defparam ii3079.CONFIG_DATA = 16'h5555;
      defparam ii3079.PLACE_LOCATION = "NONE";
      defparam ii3079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3080 ( .DX(nn3080), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2034_), .F2(dummy_abc_2035_), .F3(dummy_abc_2036_) );
      defparam ii3080.CONFIG_DATA = 16'h5555;
      defparam ii3080.PLACE_LOCATION = "NONE";
      defparam ii3080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3081 ( .DX(nn3081), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2037_), .F2(dummy_abc_2038_), .F3(dummy_abc_2039_) );
      defparam ii3081.CONFIG_DATA = 16'h5555;
      defparam ii3081.PLACE_LOCATION = "NONE";
      defparam ii3081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3082 ( .DX(nn3082), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2040_), .F2(dummy_abc_2041_), .F3(dummy_abc_2042_) );
      defparam ii3082.CONFIG_DATA = 16'h5555;
      defparam ii3082.PLACE_LOCATION = "NONE";
      defparam ii3082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3083 ( .DX(nn3083), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2043_), .F2(dummy_abc_2044_), .F3(dummy_abc_2045_) );
      defparam ii3083.CONFIG_DATA = 16'h5555;
      defparam ii3083.PLACE_LOCATION = "NONE";
      defparam ii3083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3084 ( .DX(nn3084), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2046_), .F2(dummy_abc_2047_), .F3(dummy_abc_2048_) );
      defparam ii3084.CONFIG_DATA = 16'h5555;
      defparam ii3084.PLACE_LOCATION = "NONE";
      defparam ii3084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3085 ( .DX(nn3085), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2049_), .F2(dummy_abc_2050_), .F3(dummy_abc_2051_) );
      defparam ii3085.CONFIG_DATA = 16'h5555;
      defparam ii3085.PLACE_LOCATION = "NONE";
      defparam ii3085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3086 ( .DX(nn3086), .F0(dummy_abc_2052_), .F1(dummy_abc_2053_), .F2(dummy_abc_2054_), .F3(dummy_abc_2055_) );
      defparam ii3086.CONFIG_DATA = 16'hFFFF;
      defparam ii3086.PLACE_LOCATION = "NONE";
      defparam ii3086.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_231_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_261_ ), 
        .DX( {nn3086, nn3085, nn3084, nn3083, nn3082, nn3081, nn3080, nn3079, 
              nn3078, nn3077, nn3076, nn3075, nn3074, nn3073, nn3072, nn3071, 
              nn3032, nn3031} ), 
        .SUM( {\coefcal1_divide_inst1_u124_XORCI_17|SUM_net , dummy_262_, 
              dummy_263_, dummy_264_, dummy_265_, dummy_266_, dummy_267_, dummy_268_, 
              dummy_269_, dummy_270_, dummy_271_, dummy_272_, dummy_273_, dummy_274_, 
              dummy_275_, dummy_276_, dummy_277_, dummy_278_} )
      );
    CS_LUT4_PRIM ii3107 ( .DX(nn3107), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_242_), .F3(dummy_abc_2056_) );
      defparam ii3107.CONFIG_DATA = 16'hA6A6;
      defparam ii3107.PLACE_LOCATION = "NONE";
      defparam ii3107.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3108 ( .DX(nn3108), .F0(dummy_242_), .F1(nn3033), .F2(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ), .F3(dummy_abc_2057_) );
      defparam ii3108.CONFIG_DATA = 16'hD8D8;
      defparam ii3108.PLACE_LOCATION = "NONE";
      defparam ii3108.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3109 ( .DX(nn3109), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2058_), .F3(dummy_abc_2059_) );
      defparam ii3109.CONFIG_DATA = 16'h9999;
      defparam ii3109.PLACE_LOCATION = "NONE";
      defparam ii3109.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3110 ( .DX(nn3110), .F0(\coefcal1_xDividend__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_242_) );
      defparam ii3110.CONFIG_DATA = 16'hA569;
      defparam ii3110.PLACE_LOCATION = "NONE";
      defparam ii3110.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3111 ( .DX(nn3111), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_242_), .F2(nn3033), .F3(\coefcal1_divide_inst1_u103_XORCI_1|SUM_net ) );
      defparam ii3111.CONFIG_DATA = 16'hA695;
      defparam ii3111.PLACE_LOCATION = "NONE";
      defparam ii3111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3112 ( .DX(nn3112), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3034), .F2(dummy_242_), .F3(\coefcal1_divide_inst1_u103_XORCI_2|SUM_net ) );
      defparam ii3112.CONFIG_DATA = 16'h9A95;
      defparam ii3112.PLACE_LOCATION = "NONE";
      defparam ii3112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3113 ( .DX(nn3113), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_abc_2060_), .F2(dummy_abc_2061_), .F3(dummy_abc_2062_) );
      defparam ii3113.CONFIG_DATA = 16'h5555;
      defparam ii3113.PLACE_LOCATION = "NONE";
      defparam ii3113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3114 ( .DX(nn3114), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_2063_), .F2(dummy_abc_2064_), .F3(dummy_abc_2065_) );
      defparam ii3114.CONFIG_DATA = 16'h5555;
      defparam ii3114.PLACE_LOCATION = "NONE";
      defparam ii3114.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3115 ( .DX(nn3115), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2066_), .F2(dummy_abc_2067_), .F3(dummy_abc_2068_) );
      defparam ii3115.CONFIG_DATA = 16'h5555;
      defparam ii3115.PLACE_LOCATION = "NONE";
      defparam ii3115.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3116 ( .DX(nn3116), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2069_), .F2(dummy_abc_2070_), .F3(dummy_abc_2071_) );
      defparam ii3116.CONFIG_DATA = 16'h5555;
      defparam ii3116.PLACE_LOCATION = "NONE";
      defparam ii3116.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3117 ( .DX(nn3117), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2072_), .F2(dummy_abc_2073_), .F3(dummy_abc_2074_) );
      defparam ii3117.CONFIG_DATA = 16'h5555;
      defparam ii3117.PLACE_LOCATION = "NONE";
      defparam ii3117.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3118 ( .DX(nn3118), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2075_), .F2(dummy_abc_2076_), .F3(dummy_abc_2077_) );
      defparam ii3118.CONFIG_DATA = 16'h5555;
      defparam ii3118.PLACE_LOCATION = "NONE";
      defparam ii3118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3119 ( .DX(nn3119), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2078_), .F2(dummy_abc_2079_), .F3(dummy_abc_2080_) );
      defparam ii3119.CONFIG_DATA = 16'h5555;
      defparam ii3119.PLACE_LOCATION = "NONE";
      defparam ii3119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3120 ( .DX(nn3120), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2081_), .F2(dummy_abc_2082_), .F3(dummy_abc_2083_) );
      defparam ii3120.CONFIG_DATA = 16'h5555;
      defparam ii3120.PLACE_LOCATION = "NONE";
      defparam ii3120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3121 ( .DX(nn3121), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2084_), .F2(dummy_abc_2085_), .F3(dummy_abc_2086_) );
      defparam ii3121.CONFIG_DATA = 16'h5555;
      defparam ii3121.PLACE_LOCATION = "NONE";
      defparam ii3121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3122 ( .DX(nn3122), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2087_), .F2(dummy_abc_2088_), .F3(dummy_abc_2089_) );
      defparam ii3122.CONFIG_DATA = 16'h5555;
      defparam ii3122.PLACE_LOCATION = "NONE";
      defparam ii3122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3123 ( .DX(nn3123), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2090_), .F2(dummy_abc_2091_), .F3(dummy_abc_2092_) );
      defparam ii3123.CONFIG_DATA = 16'h5555;
      defparam ii3123.PLACE_LOCATION = "NONE";
      defparam ii3123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3124 ( .DX(nn3124), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2093_), .F2(dummy_abc_2094_), .F3(dummy_abc_2095_) );
      defparam ii3124.CONFIG_DATA = 16'h5555;
      defparam ii3124.PLACE_LOCATION = "NONE";
      defparam ii3124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3125 ( .DX(nn3125), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2096_), .F2(dummy_abc_2097_), .F3(dummy_abc_2098_) );
      defparam ii3125.CONFIG_DATA = 16'h5555;
      defparam ii3125.PLACE_LOCATION = "NONE";
      defparam ii3125.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_216_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3108, 
              nn3107, \coefcal1_xDividend__reg[13]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_145_ ), 
        .DX( {nn3125, nn3124, nn3123, nn3122, nn3121, nn3120, nn3119, nn3118, 
              nn3117, nn3116, nn3115, nn3114, nn3113, nn3112, nn3111, nn3110, 
              nn3109} ), 
        .SUM( {dummy_146_, \coefcal1_divide_inst1_u104_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_14|SUM_net , \coefcal1_divide_inst1_u104_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_12|SUM_net , \coefcal1_divide_inst1_u104_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_10|SUM_net , \coefcal1_divide_inst1_u104_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_8|SUM_net , \coefcal1_divide_inst1_u104_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_6|SUM_net , \coefcal1_divide_inst1_u104_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_4|SUM_net , \coefcal1_divide_inst1_u104_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_2|SUM_net , \coefcal1_divide_inst1_u104_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u104_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3145 ( .DX(nn3145), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(dummy_242_), .F2(dummy_261_), .F3(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ) );
      defparam ii3145.CONFIG_DATA = 16'h8A80;
      defparam ii3145.PLACE_LOCATION = "NONE";
      defparam ii3145.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3146 ( .DX(nn3146), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2099_), .F3(dummy_abc_2100_) );
      defparam ii3146.CONFIG_DATA = 16'h9999;
      defparam ii3146.PLACE_LOCATION = "NONE";
      defparam ii3146.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3147 ( .DX(nn3147), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_261_) );
      defparam ii3147.CONFIG_DATA = 16'hA569;
      defparam ii3147.PLACE_LOCATION = "NONE";
      defparam ii3147.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3148 ( .DX(nn3148), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_261_), .F2(nn3107), .F3(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ) );
      defparam ii3148.CONFIG_DATA = 16'hA695;
      defparam ii3148.PLACE_LOCATION = "NONE";
      defparam ii3148.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3149 ( .DX(nn3149), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3108), .F2(dummy_261_), .F3(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ) );
      defparam ii3149.CONFIG_DATA = 16'h9A95;
      defparam ii3149.PLACE_LOCATION = "NONE";
      defparam ii3149.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3150 ( .DX(nn3150), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(dummy_242_), .F2(dummy_261_), .F3(dummy_abc_2101_) );
      defparam ii3150.CONFIG_DATA = 16'h8A8A;
      defparam ii3150.PLACE_LOCATION = "NONE";
      defparam ii3150.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3151 ( .DX(nn3151), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_261_), .F2(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ), .F3(nn3150) );
      defparam ii3151.CONFIG_DATA = 16'hA955;
      defparam ii3151.PLACE_LOCATION = "NONE";
      defparam ii3151.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3152 ( .DX(nn3152), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_2102_), .F2(dummy_abc_2103_), .F3(dummy_abc_2104_) );
      defparam ii3152.CONFIG_DATA = 16'h5555;
      defparam ii3152.PLACE_LOCATION = "NONE";
      defparam ii3152.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3153 ( .DX(nn3153), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2105_), .F2(dummy_abc_2106_), .F3(dummy_abc_2107_) );
      defparam ii3153.CONFIG_DATA = 16'h5555;
      defparam ii3153.PLACE_LOCATION = "NONE";
      defparam ii3153.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3154 ( .DX(nn3154), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2108_), .F2(dummy_abc_2109_), .F3(dummy_abc_2110_) );
      defparam ii3154.CONFIG_DATA = 16'h5555;
      defparam ii3154.PLACE_LOCATION = "NONE";
      defparam ii3154.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3155 ( .DX(nn3155), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2111_), .F2(dummy_abc_2112_), .F3(dummy_abc_2113_) );
      defparam ii3155.CONFIG_DATA = 16'h5555;
      defparam ii3155.PLACE_LOCATION = "NONE";
      defparam ii3155.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3156 ( .DX(nn3156), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2114_), .F2(dummy_abc_2115_), .F3(dummy_abc_2116_) );
      defparam ii3156.CONFIG_DATA = 16'h5555;
      defparam ii3156.PLACE_LOCATION = "NONE";
      defparam ii3156.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3157 ( .DX(nn3157), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2117_), .F2(dummy_abc_2118_), .F3(dummy_abc_2119_) );
      defparam ii3157.CONFIG_DATA = 16'h5555;
      defparam ii3157.PLACE_LOCATION = "NONE";
      defparam ii3157.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3158 ( .DX(nn3158), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2120_), .F2(dummy_abc_2121_), .F3(dummy_abc_2122_) );
      defparam ii3158.CONFIG_DATA = 16'h5555;
      defparam ii3158.PLACE_LOCATION = "NONE";
      defparam ii3158.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3159 ( .DX(nn3159), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2123_), .F2(dummy_abc_2124_), .F3(dummy_abc_2125_) );
      defparam ii3159.CONFIG_DATA = 16'h5555;
      defparam ii3159.PLACE_LOCATION = "NONE";
      defparam ii3159.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3160 ( .DX(nn3160), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2126_), .F2(dummy_abc_2127_), .F3(dummy_abc_2128_) );
      defparam ii3160.CONFIG_DATA = 16'h5555;
      defparam ii3160.PLACE_LOCATION = "NONE";
      defparam ii3160.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3161 ( .DX(nn3161), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2129_), .F2(dummy_abc_2130_), .F3(dummy_abc_2131_) );
      defparam ii3161.CONFIG_DATA = 16'h5555;
      defparam ii3161.PLACE_LOCATION = "NONE";
      defparam ii3161.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3162 ( .DX(nn3162), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2132_), .F2(dummy_abc_2133_), .F3(dummy_abc_2134_) );
      defparam ii3162.CONFIG_DATA = 16'h5555;
      defparam ii3162.PLACE_LOCATION = "NONE";
      defparam ii3162.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3163 ( .DX(nn3163), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2135_), .F2(dummy_abc_2136_), .F3(dummy_abc_2137_) );
      defparam ii3163.CONFIG_DATA = 16'h5555;
      defparam ii3163.PLACE_LOCATION = "NONE";
      defparam ii3163.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3164 ( .DX(nn3164), .F0(dummy_abc_2138_), .F1(dummy_abc_2139_), .F2(dummy_abc_2140_), .F3(dummy_abc_2141_) );
      defparam ii3164.CONFIG_DATA = 16'hFFFF;
      defparam ii3164.PLACE_LOCATION = "NONE";
      defparam ii3164.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_232_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_280_ ), 
        .DX( {nn3164, nn3163, nn3162, nn3161, nn3160, nn3159, nn3158, nn3157, 
              nn3156, nn3155, nn3154, nn3153, nn3152, nn3151, nn3149, nn3148, 
              nn3147, nn3146} ), 
        .SUM( {\coefcal1_divide_inst1_u126_XORCI_17|SUM_net , dummy_281_, 
              dummy_282_, dummy_283_, dummy_284_, dummy_285_, dummy_286_, dummy_287_, 
              dummy_288_, dummy_289_, dummy_290_, dummy_291_, dummy_292_, dummy_293_, 
              dummy_294_, dummy_295_, dummy_296_, dummy_297_} )
      );
    CS_LUT4_PRIM ii3185 ( .DX(nn3185), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2142_), .F3(dummy_abc_2143_) );
      defparam ii3185.CONFIG_DATA = 16'h9999;
      defparam ii3185.PLACE_LOCATION = "NONE";
      defparam ii3185.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3186 ( .DX(nn3186), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_280_) );
      defparam ii3186.CONFIG_DATA = 16'hA569;
      defparam ii3186.PLACE_LOCATION = "NONE";
      defparam ii3186.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3187 ( .DX(nn3187), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_261_), .F3(dummy_abc_2144_) );
      defparam ii3187.CONFIG_DATA = 16'hA6A6;
      defparam ii3187.PLACE_LOCATION = "NONE";
      defparam ii3187.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3188 ( .DX(nn3188), .F0(dummy_261_), .F1(nn3107), .F2(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ), .F3(dummy_abc_2145_) );
      defparam ii3188.CONFIG_DATA = 16'hD8D8;
      defparam ii3188.PLACE_LOCATION = "NONE";
      defparam ii3188.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3189 ( .DX(nn3189), .F0(nn3108), .F1(dummy_261_), .F2(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ), .F3(dummy_abc_2146_) );
      defparam ii3189.CONFIG_DATA = 16'hB8B8;
      defparam ii3189.PLACE_LOCATION = "NONE";
      defparam ii3189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3190 ( .DX(nn3190), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2147_), .F3(dummy_abc_2148_) );
      defparam ii3190.CONFIG_DATA = 16'h9999;
      defparam ii3190.PLACE_LOCATION = "NONE";
      defparam ii3190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3191 ( .DX(nn3191), .F0(\coefcal1_xDividend__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_261_) );
      defparam ii3191.CONFIG_DATA = 16'hA569;
      defparam ii3191.PLACE_LOCATION = "NONE";
      defparam ii3191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3192 ( .DX(nn3192), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_261_), .F2(nn3107), .F3(\coefcal1_divide_inst1_u104_XORCI_1|SUM_net ) );
      defparam ii3192.CONFIG_DATA = 16'hA695;
      defparam ii3192.PLACE_LOCATION = "NONE";
      defparam ii3192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3193 ( .DX(nn3193), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3108), .F2(dummy_261_), .F3(\coefcal1_divide_inst1_u104_XORCI_2|SUM_net ) );
      defparam ii3193.CONFIG_DATA = 16'h9A95;
      defparam ii3193.PLACE_LOCATION = "NONE";
      defparam ii3193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3194 ( .DX(nn3194), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(dummy_261_), .F2(\coefcal1_divide_inst1_u104_XORCI_3|SUM_net ), .F3(nn3150) );
      defparam ii3194.CONFIG_DATA = 16'hA955;
      defparam ii3194.PLACE_LOCATION = "NONE";
      defparam ii3194.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3195 ( .DX(nn3195), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(dummy_abc_2149_), .F2(dummy_abc_2150_), .F3(dummy_abc_2151_) );
      defparam ii3195.CONFIG_DATA = 16'h5555;
      defparam ii3195.PLACE_LOCATION = "NONE";
      defparam ii3195.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3196 ( .DX(nn3196), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2152_), .F2(dummy_abc_2153_), .F3(dummy_abc_2154_) );
      defparam ii3196.CONFIG_DATA = 16'h5555;
      defparam ii3196.PLACE_LOCATION = "NONE";
      defparam ii3196.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3197 ( .DX(nn3197), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2155_), .F2(dummy_abc_2156_), .F3(dummy_abc_2157_) );
      defparam ii3197.CONFIG_DATA = 16'h5555;
      defparam ii3197.PLACE_LOCATION = "NONE";
      defparam ii3197.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3198 ( .DX(nn3198), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2158_), .F2(dummy_abc_2159_), .F3(dummy_abc_2160_) );
      defparam ii3198.CONFIG_DATA = 16'h5555;
      defparam ii3198.PLACE_LOCATION = "NONE";
      defparam ii3198.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3199 ( .DX(nn3199), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2161_), .F2(dummy_abc_2162_), .F3(dummy_abc_2163_) );
      defparam ii3199.CONFIG_DATA = 16'h5555;
      defparam ii3199.PLACE_LOCATION = "NONE";
      defparam ii3199.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3200 ( .DX(nn3200), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2164_), .F2(dummy_abc_2165_), .F3(dummy_abc_2166_) );
      defparam ii3200.CONFIG_DATA = 16'h5555;
      defparam ii3200.PLACE_LOCATION = "NONE";
      defparam ii3200.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3201 ( .DX(nn3201), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2167_), .F2(dummy_abc_2168_), .F3(dummy_abc_2169_) );
      defparam ii3201.CONFIG_DATA = 16'h5555;
      defparam ii3201.PLACE_LOCATION = "NONE";
      defparam ii3201.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3202 ( .DX(nn3202), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2170_), .F2(dummy_abc_2171_), .F3(dummy_abc_2172_) );
      defparam ii3202.CONFIG_DATA = 16'h5555;
      defparam ii3202.PLACE_LOCATION = "NONE";
      defparam ii3202.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3203 ( .DX(nn3203), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2173_), .F2(dummy_abc_2174_), .F3(dummy_abc_2175_) );
      defparam ii3203.CONFIG_DATA = 16'h5555;
      defparam ii3203.PLACE_LOCATION = "NONE";
      defparam ii3203.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3204 ( .DX(nn3204), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2176_), .F2(dummy_abc_2177_), .F3(dummy_abc_2178_) );
      defparam ii3204.CONFIG_DATA = 16'h5555;
      defparam ii3204.PLACE_LOCATION = "NONE";
      defparam ii3204.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3205 ( .DX(nn3205), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2179_), .F2(dummy_abc_2180_), .F3(dummy_abc_2181_) );
      defparam ii3205.CONFIG_DATA = 16'h5555;
      defparam ii3205.PLACE_LOCATION = "NONE";
      defparam ii3205.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3206 ( .DX(nn3206), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2182_), .F2(dummy_abc_2183_), .F3(dummy_abc_2184_) );
      defparam ii3206.CONFIG_DATA = 16'h5555;
      defparam ii3206.PLACE_LOCATION = "NONE";
      defparam ii3206.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_217_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn3145, nn3189, nn3188, nn3187, 
              \coefcal1_xDividend__reg[12]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_147_ ), 
        .DX( {nn3206, nn3205, nn3204, nn3203, nn3202, nn3201, nn3200, nn3199, 
              nn3198, nn3197, nn3196, nn3195, nn3194, nn3193, nn3192, nn3191, 
              nn3190} ), 
        .SUM( {dummy_148_, \coefcal1_divide_inst1_u105_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_14|SUM_net , \coefcal1_divide_inst1_u105_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_12|SUM_net , \coefcal1_divide_inst1_u105_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_10|SUM_net , \coefcal1_divide_inst1_u105_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_8|SUM_net , \coefcal1_divide_inst1_u105_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_6|SUM_net , \coefcal1_divide_inst1_u105_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_4|SUM_net , \coefcal1_divide_inst1_u105_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_2|SUM_net , \coefcal1_divide_inst1_u105_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u105_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3226 ( .DX(nn3226), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_280_), .F2(nn3187), .F3(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ) );
      defparam ii3226.CONFIG_DATA = 16'hA695;
      defparam ii3226.PLACE_LOCATION = "NONE";
      defparam ii3226.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3227 ( .DX(nn3227), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3188), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ) );
      defparam ii3227.CONFIG_DATA = 16'h9A95;
      defparam ii3227.PLACE_LOCATION = "NONE";
      defparam ii3227.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3228 ( .DX(nn3228), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3189), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ) );
      defparam ii3228.CONFIG_DATA = 16'h9A95;
      defparam ii3228.PLACE_LOCATION = "NONE";
      defparam ii3228.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3229 ( .DX(nn3229), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3145), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_4|SUM_net ) );
      defparam ii3229.CONFIG_DATA = 16'h9A95;
      defparam ii3229.PLACE_LOCATION = "NONE";
      defparam ii3229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3230 ( .DX(nn3230), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2185_), .F2(dummy_abc_2186_), .F3(dummy_abc_2187_) );
      defparam ii3230.CONFIG_DATA = 16'h5555;
      defparam ii3230.PLACE_LOCATION = "NONE";
      defparam ii3230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3231 ( .DX(nn3231), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2188_), .F2(dummy_abc_2189_), .F3(dummy_abc_2190_) );
      defparam ii3231.CONFIG_DATA = 16'h5555;
      defparam ii3231.PLACE_LOCATION = "NONE";
      defparam ii3231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3232 ( .DX(nn3232), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2191_), .F2(dummy_abc_2192_), .F3(dummy_abc_2193_) );
      defparam ii3232.CONFIG_DATA = 16'h5555;
      defparam ii3232.PLACE_LOCATION = "NONE";
      defparam ii3232.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3233 ( .DX(nn3233), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2194_), .F2(dummy_abc_2195_), .F3(dummy_abc_2196_) );
      defparam ii3233.CONFIG_DATA = 16'h5555;
      defparam ii3233.PLACE_LOCATION = "NONE";
      defparam ii3233.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3234 ( .DX(nn3234), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2197_), .F2(dummy_abc_2198_), .F3(dummy_abc_2199_) );
      defparam ii3234.CONFIG_DATA = 16'h5555;
      defparam ii3234.PLACE_LOCATION = "NONE";
      defparam ii3234.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3235 ( .DX(nn3235), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2200_), .F2(dummy_abc_2201_), .F3(dummy_abc_2202_) );
      defparam ii3235.CONFIG_DATA = 16'h5555;
      defparam ii3235.PLACE_LOCATION = "NONE";
      defparam ii3235.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3236 ( .DX(nn3236), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2203_), .F2(dummy_abc_2204_), .F3(dummy_abc_2205_) );
      defparam ii3236.CONFIG_DATA = 16'h5555;
      defparam ii3236.PLACE_LOCATION = "NONE";
      defparam ii3236.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3237 ( .DX(nn3237), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2206_), .F2(dummy_abc_2207_), .F3(dummy_abc_2208_) );
      defparam ii3237.CONFIG_DATA = 16'h5555;
      defparam ii3237.PLACE_LOCATION = "NONE";
      defparam ii3237.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3238 ( .DX(nn3238), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2209_), .F2(dummy_abc_2210_), .F3(dummy_abc_2211_) );
      defparam ii3238.CONFIG_DATA = 16'h5555;
      defparam ii3238.PLACE_LOCATION = "NONE";
      defparam ii3238.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3239 ( .DX(nn3239), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2212_), .F2(dummy_abc_2213_), .F3(dummy_abc_2214_) );
      defparam ii3239.CONFIG_DATA = 16'h5555;
      defparam ii3239.PLACE_LOCATION = "NONE";
      defparam ii3239.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3240 ( .DX(nn3240), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2215_), .F2(dummy_abc_2216_), .F3(dummy_abc_2217_) );
      defparam ii3240.CONFIG_DATA = 16'h5555;
      defparam ii3240.PLACE_LOCATION = "NONE";
      defparam ii3240.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3241 ( .DX(nn3241), .F0(dummy_abc_2218_), .F1(dummy_abc_2219_), .F2(dummy_abc_2220_), .F3(dummy_abc_2221_) );
      defparam ii3241.CONFIG_DATA = 16'hFFFF;
      defparam ii3241.PLACE_LOCATION = "NONE";
      defparam ii3241.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_233_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_299_ ), 
        .DX( {nn3241, nn3240, nn3239, nn3238, nn3237, nn3236, nn3235, nn3234, 
              nn3233, nn3232, nn3231, nn3230, nn3229, nn3228, nn3227, nn3226, 
              nn3186, nn3185} ), 
        .SUM( {\coefcal1_divide_inst1_u128_XORCI_17|SUM_net , dummy_300_, 
              dummy_301_, dummy_302_, dummy_303_, dummy_304_, dummy_305_, dummy_306_, 
              dummy_307_, dummy_308_, dummy_309_, dummy_310_, dummy_311_, dummy_312_, 
              dummy_313_, dummy_314_, dummy_315_, dummy_316_} )
      );
    CS_LUT4_PRIM ii3262 ( .DX(nn3262), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_280_), .F3(dummy_abc_2222_) );
      defparam ii3262.CONFIG_DATA = 16'hA6A6;
      defparam ii3262.PLACE_LOCATION = "NONE";
      defparam ii3262.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3263 ( .DX(nn3263), .F0(dummy_280_), .F1(nn3187), .F2(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ), .F3(dummy_abc_2223_) );
      defparam ii3263.CONFIG_DATA = 16'hD8D8;
      defparam ii3263.PLACE_LOCATION = "NONE";
      defparam ii3263.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3264 ( .DX(nn3264), .F0(nn3188), .F1(dummy_280_), .F2(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ), .F3(dummy_abc_2224_) );
      defparam ii3264.CONFIG_DATA = 16'hB8B8;
      defparam ii3264.PLACE_LOCATION = "NONE";
      defparam ii3264.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3265 ( .DX(nn3265), .F0(nn3189), .F1(dummy_280_), .F2(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ), .F3(dummy_abc_2225_) );
      defparam ii3265.CONFIG_DATA = 16'hB8B8;
      defparam ii3265.PLACE_LOCATION = "NONE";
      defparam ii3265.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3266 ( .DX(nn3266), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2226_), .F3(dummy_abc_2227_) );
      defparam ii3266.CONFIG_DATA = 16'h9999;
      defparam ii3266.PLACE_LOCATION = "NONE";
      defparam ii3266.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3267 ( .DX(nn3267), .F0(\coefcal1_xDividend__reg[12]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_280_) );
      defparam ii3267.CONFIG_DATA = 16'hA569;
      defparam ii3267.PLACE_LOCATION = "NONE";
      defparam ii3267.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3268 ( .DX(nn3268), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_280_), .F2(nn3187), .F3(\coefcal1_divide_inst1_u105_XORCI_1|SUM_net ) );
      defparam ii3268.CONFIG_DATA = 16'hA695;
      defparam ii3268.PLACE_LOCATION = "NONE";
      defparam ii3268.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3269 ( .DX(nn3269), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3188), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_2|SUM_net ) );
      defparam ii3269.CONFIG_DATA = 16'h9A95;
      defparam ii3269.PLACE_LOCATION = "NONE";
      defparam ii3269.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3270 ( .DX(nn3270), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3189), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_3|SUM_net ) );
      defparam ii3270.CONFIG_DATA = 16'h9A95;
      defparam ii3270.PLACE_LOCATION = "NONE";
      defparam ii3270.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3271 ( .DX(nn3271), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3145), .F2(dummy_280_), .F3(\coefcal1_divide_inst1_u105_XORCI_4|SUM_net ) );
      defparam ii3271.CONFIG_DATA = 16'h9A95;
      defparam ii3271.PLACE_LOCATION = "NONE";
      defparam ii3271.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3272 ( .DX(nn3272), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(dummy_abc_2228_), .F2(dummy_abc_2229_), .F3(dummy_abc_2230_) );
      defparam ii3272.CONFIG_DATA = 16'h5555;
      defparam ii3272.PLACE_LOCATION = "NONE";
      defparam ii3272.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3273 ( .DX(nn3273), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2231_), .F2(dummy_abc_2232_), .F3(dummy_abc_2233_) );
      defparam ii3273.CONFIG_DATA = 16'h5555;
      defparam ii3273.PLACE_LOCATION = "NONE";
      defparam ii3273.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3274 ( .DX(nn3274), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2234_), .F2(dummy_abc_2235_), .F3(dummy_abc_2236_) );
      defparam ii3274.CONFIG_DATA = 16'h5555;
      defparam ii3274.PLACE_LOCATION = "NONE";
      defparam ii3274.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3275 ( .DX(nn3275), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2237_), .F2(dummy_abc_2238_), .F3(dummy_abc_2239_) );
      defparam ii3275.CONFIG_DATA = 16'h5555;
      defparam ii3275.PLACE_LOCATION = "NONE";
      defparam ii3275.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3276 ( .DX(nn3276), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2240_), .F2(dummy_abc_2241_), .F3(dummy_abc_2242_) );
      defparam ii3276.CONFIG_DATA = 16'h5555;
      defparam ii3276.PLACE_LOCATION = "NONE";
      defparam ii3276.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3277 ( .DX(nn3277), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2243_), .F2(dummy_abc_2244_), .F3(dummy_abc_2245_) );
      defparam ii3277.CONFIG_DATA = 16'h5555;
      defparam ii3277.PLACE_LOCATION = "NONE";
      defparam ii3277.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3278 ( .DX(nn3278), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2246_), .F2(dummy_abc_2247_), .F3(dummy_abc_2248_) );
      defparam ii3278.CONFIG_DATA = 16'h5555;
      defparam ii3278.PLACE_LOCATION = "NONE";
      defparam ii3278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3279 ( .DX(nn3279), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2249_), .F2(dummy_abc_2250_), .F3(dummy_abc_2251_) );
      defparam ii3279.CONFIG_DATA = 16'h5555;
      defparam ii3279.PLACE_LOCATION = "NONE";
      defparam ii3279.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3280 ( .DX(nn3280), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2252_), .F2(dummy_abc_2253_), .F3(dummy_abc_2254_) );
      defparam ii3280.CONFIG_DATA = 16'h5555;
      defparam ii3280.PLACE_LOCATION = "NONE";
      defparam ii3280.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3281 ( .DX(nn3281), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2255_), .F2(dummy_abc_2256_), .F3(dummy_abc_2257_) );
      defparam ii3281.CONFIG_DATA = 16'h5555;
      defparam ii3281.PLACE_LOCATION = "NONE";
      defparam ii3281.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3282 ( .DX(nn3282), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2258_), .F2(dummy_abc_2259_), .F3(dummy_abc_2260_) );
      defparam ii3282.CONFIG_DATA = 16'h5555;
      defparam ii3282.PLACE_LOCATION = "NONE";
      defparam ii3282.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_218_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn3265, nn3264, nn3263, nn3262, 
              \coefcal1_xDividend__reg[11]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_149_ ), 
        .DX( {nn3282, nn3281, nn3280, nn3279, nn3278, nn3277, nn3276, nn3275, 
              nn3274, nn3273, nn3272, nn3271, nn3270, nn3269, nn3268, nn3267, 
              nn3266} ), 
        .SUM( {dummy_150_, \coefcal1_divide_inst1_u106_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_14|SUM_net , \coefcal1_divide_inst1_u106_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_12|SUM_net , \coefcal1_divide_inst1_u106_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_10|SUM_net , \coefcal1_divide_inst1_u106_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_8|SUM_net , \coefcal1_divide_inst1_u106_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_6|SUM_net , \coefcal1_divide_inst1_u106_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_4|SUM_net , \coefcal1_divide_inst1_u106_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_2|SUM_net , \coefcal1_divide_inst1_u106_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u106_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3302 ( .DX(nn3302), .F0(nn3145), .F1(dummy_280_), .F2(dummy_299_), .F3(\coefcal1_divide_inst1_u106_XORCI_5|SUM_net ) );
      defparam ii3302.CONFIG_DATA = 16'h8A80;
      defparam ii3302.PLACE_LOCATION = "NONE";
      defparam ii3302.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3303 ( .DX(nn3303), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2261_), .F3(dummy_abc_2262_) );
      defparam ii3303.CONFIG_DATA = 16'h9999;
      defparam ii3303.PLACE_LOCATION = "NONE";
      defparam ii3303.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3304 ( .DX(nn3304), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_299_) );
      defparam ii3304.CONFIG_DATA = 16'hA569;
      defparam ii3304.PLACE_LOCATION = "NONE";
      defparam ii3304.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3305 ( .DX(nn3305), .F0(dummy_299_), .F1(nn3262), .F2(\coefcal1_divide_inst1_u106_XORCI_1|SUM_net ), .F3(dummy_abc_2263_) );
      defparam ii3305.CONFIG_DATA = 16'hD8D8;
      defparam ii3305.PLACE_LOCATION = "NONE";
      defparam ii3305.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3306 ( .DX(nn3306), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(nn3305), .F2(dummy_abc_2264_), .F3(dummy_abc_2265_) );
      defparam ii3306.CONFIG_DATA = 16'h9999;
      defparam ii3306.PLACE_LOCATION = "NONE";
      defparam ii3306.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3307 ( .DX(nn3307), .F0(nn3263), .F1(dummy_299_), .F2(\coefcal1_divide_inst1_u106_XORCI_2|SUM_net ), .F3(dummy_abc_2266_) );
      defparam ii3307.CONFIG_DATA = 16'hB8B8;
      defparam ii3307.PLACE_LOCATION = "NONE";
      defparam ii3307.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3308 ( .DX(nn3308), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3307), .F2(dummy_abc_2267_), .F3(dummy_abc_2268_) );
      defparam ii3308.CONFIG_DATA = 16'h9999;
      defparam ii3308.PLACE_LOCATION = "NONE";
      defparam ii3308.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3309 ( .DX(nn3309), .F0(nn3264), .F1(dummy_299_), .F2(\coefcal1_divide_inst1_u106_XORCI_3|SUM_net ), .F3(dummy_abc_2269_) );
      defparam ii3309.CONFIG_DATA = 16'hB8B8;
      defparam ii3309.PLACE_LOCATION = "NONE";
      defparam ii3309.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3310 ( .DX(nn3310), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3309), .F2(dummy_abc_2270_), .F3(dummy_abc_2271_) );
      defparam ii3310.CONFIG_DATA = 16'h9999;
      defparam ii3310.PLACE_LOCATION = "NONE";
      defparam ii3310.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3311 ( .DX(nn3311), .F0(nn3265), .F1(dummy_299_), .F2(\coefcal1_divide_inst1_u106_XORCI_4|SUM_net ), .F3(dummy_abc_2272_) );
      defparam ii3311.CONFIG_DATA = 16'hB8B8;
      defparam ii3311.PLACE_LOCATION = "NONE";
      defparam ii3311.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3312 ( .DX(nn3312), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3311), .F2(dummy_abc_2273_), .F3(dummy_abc_2274_) );
      defparam ii3312.CONFIG_DATA = 16'h9999;
      defparam ii3312.PLACE_LOCATION = "NONE";
      defparam ii3312.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3313 ( .DX(nn3313), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3302), .F2(dummy_abc_2275_), .F3(dummy_abc_2276_) );
      defparam ii3313.CONFIG_DATA = 16'h9999;
      defparam ii3313.PLACE_LOCATION = "NONE";
      defparam ii3313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3314 ( .DX(nn3314), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2277_), .F2(dummy_abc_2278_), .F3(dummy_abc_2279_) );
      defparam ii3314.CONFIG_DATA = 16'h5555;
      defparam ii3314.PLACE_LOCATION = "NONE";
      defparam ii3314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3315 ( .DX(nn3315), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2280_), .F2(dummy_abc_2281_), .F3(dummy_abc_2282_) );
      defparam ii3315.CONFIG_DATA = 16'h5555;
      defparam ii3315.PLACE_LOCATION = "NONE";
      defparam ii3315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3316 ( .DX(nn3316), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2283_), .F2(dummy_abc_2284_), .F3(dummy_abc_2285_) );
      defparam ii3316.CONFIG_DATA = 16'h5555;
      defparam ii3316.PLACE_LOCATION = "NONE";
      defparam ii3316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3317 ( .DX(nn3317), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2286_), .F2(dummy_abc_2287_), .F3(dummy_abc_2288_) );
      defparam ii3317.CONFIG_DATA = 16'h5555;
      defparam ii3317.PLACE_LOCATION = "NONE";
      defparam ii3317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3318 ( .DX(nn3318), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2289_), .F2(dummy_abc_2290_), .F3(dummy_abc_2291_) );
      defparam ii3318.CONFIG_DATA = 16'h5555;
      defparam ii3318.PLACE_LOCATION = "NONE";
      defparam ii3318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3319 ( .DX(nn3319), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2292_), .F2(dummy_abc_2293_), .F3(dummy_abc_2294_) );
      defparam ii3319.CONFIG_DATA = 16'h5555;
      defparam ii3319.PLACE_LOCATION = "NONE";
      defparam ii3319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3320 ( .DX(nn3320), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2295_), .F2(dummy_abc_2296_), .F3(dummy_abc_2297_) );
      defparam ii3320.CONFIG_DATA = 16'h5555;
      defparam ii3320.PLACE_LOCATION = "NONE";
      defparam ii3320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3321 ( .DX(nn3321), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2298_), .F2(dummy_abc_2299_), .F3(dummy_abc_2300_) );
      defparam ii3321.CONFIG_DATA = 16'h5555;
      defparam ii3321.PLACE_LOCATION = "NONE";
      defparam ii3321.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3322 ( .DX(nn3322), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2301_), .F2(dummy_abc_2302_), .F3(dummy_abc_2303_) );
      defparam ii3322.CONFIG_DATA = 16'h5555;
      defparam ii3322.PLACE_LOCATION = "NONE";
      defparam ii3322.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3323 ( .DX(nn3323), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2304_), .F2(dummy_abc_2305_), .F3(dummy_abc_2306_) );
      defparam ii3323.CONFIG_DATA = 16'h5555;
      defparam ii3323.PLACE_LOCATION = "NONE";
      defparam ii3323.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3324 ( .DX(nn3324), .F0(dummy_abc_2307_), .F1(dummy_abc_2308_), .F2(dummy_abc_2309_), .F3(dummy_abc_2310_) );
      defparam ii3324.CONFIG_DATA = 16'hFFFF;
      defparam ii3324.PLACE_LOCATION = "NONE";
      defparam ii3324.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_234_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_318_ ), 
        .DX( {nn3324, nn3323, nn3322, nn3321, nn3320, nn3319, nn3318, nn3317, 
              nn3316, nn3315, nn3314, nn3313, nn3312, nn3310, nn3308, nn3306, 
              nn3304, nn3303} ), 
        .SUM( {\coefcal1_divide_inst1_u130_XORCI_17|SUM_net , dummy_319_, 
              dummy_320_, dummy_321_, dummy_322_, dummy_323_, dummy_324_, dummy_325_, 
              dummy_326_, dummy_327_, dummy_328_, dummy_329_, dummy_330_, dummy_331_, 
              dummy_332_, dummy_333_, dummy_334_, dummy_335_} )
      );
    CS_LUT4_PRIM ii3345 ( .DX(nn3345), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2311_), .F3(dummy_abc_2312_) );
      defparam ii3345.CONFIG_DATA = 16'h9999;
      defparam ii3345.PLACE_LOCATION = "NONE";
      defparam ii3345.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3346 ( .DX(nn3346), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_318_) );
      defparam ii3346.CONFIG_DATA = 16'hA569;
      defparam ii3346.PLACE_LOCATION = "NONE";
      defparam ii3346.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3347 ( .DX(nn3347), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_299_), .F3(dummy_abc_2313_) );
      defparam ii3347.CONFIG_DATA = 16'hA6A6;
      defparam ii3347.PLACE_LOCATION = "NONE";
      defparam ii3347.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3348 ( .DX(nn3348), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2314_), .F3(dummy_abc_2315_) );
      defparam ii3348.CONFIG_DATA = 16'h9999;
      defparam ii3348.PLACE_LOCATION = "NONE";
      defparam ii3348.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3349 ( .DX(nn3349), .F0(\coefcal1_xDividend__reg[11]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_299_) );
      defparam ii3349.CONFIG_DATA = 16'hA569;
      defparam ii3349.PLACE_LOCATION = "NONE";
      defparam ii3349.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3350 ( .DX(nn3350), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(nn3305), .F2(dummy_abc_2316_), .F3(dummy_abc_2317_) );
      defparam ii3350.CONFIG_DATA = 16'h9999;
      defparam ii3350.PLACE_LOCATION = "NONE";
      defparam ii3350.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3351 ( .DX(nn3351), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3307), .F2(dummy_abc_2318_), .F3(dummy_abc_2319_) );
      defparam ii3351.CONFIG_DATA = 16'h9999;
      defparam ii3351.PLACE_LOCATION = "NONE";
      defparam ii3351.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3352 ( .DX(nn3352), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3309), .F2(dummy_abc_2320_), .F3(dummy_abc_2321_) );
      defparam ii3352.CONFIG_DATA = 16'h9999;
      defparam ii3352.PLACE_LOCATION = "NONE";
      defparam ii3352.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3353 ( .DX(nn3353), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3311), .F2(dummy_abc_2322_), .F3(dummy_abc_2323_) );
      defparam ii3353.CONFIG_DATA = 16'h9999;
      defparam ii3353.PLACE_LOCATION = "NONE";
      defparam ii3353.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3354 ( .DX(nn3354), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3302), .F2(dummy_abc_2324_), .F3(dummy_abc_2325_) );
      defparam ii3354.CONFIG_DATA = 16'h9999;
      defparam ii3354.PLACE_LOCATION = "NONE";
      defparam ii3354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3355 ( .DX(nn3355), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(dummy_abc_2326_), .F2(dummy_abc_2327_), .F3(dummy_abc_2328_) );
      defparam ii3355.CONFIG_DATA = 16'h5555;
      defparam ii3355.PLACE_LOCATION = "NONE";
      defparam ii3355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3356 ( .DX(nn3356), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2329_), .F2(dummy_abc_2330_), .F3(dummy_abc_2331_) );
      defparam ii3356.CONFIG_DATA = 16'h5555;
      defparam ii3356.PLACE_LOCATION = "NONE";
      defparam ii3356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3357 ( .DX(nn3357), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2332_), .F2(dummy_abc_2333_), .F3(dummy_abc_2334_) );
      defparam ii3357.CONFIG_DATA = 16'h5555;
      defparam ii3357.PLACE_LOCATION = "NONE";
      defparam ii3357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3358 ( .DX(nn3358), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2335_), .F2(dummy_abc_2336_), .F3(dummy_abc_2337_) );
      defparam ii3358.CONFIG_DATA = 16'h5555;
      defparam ii3358.PLACE_LOCATION = "NONE";
      defparam ii3358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3359 ( .DX(nn3359), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2338_), .F2(dummy_abc_2339_), .F3(dummy_abc_2340_) );
      defparam ii3359.CONFIG_DATA = 16'h5555;
      defparam ii3359.PLACE_LOCATION = "NONE";
      defparam ii3359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3360 ( .DX(nn3360), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2341_), .F2(dummy_abc_2342_), .F3(dummy_abc_2343_) );
      defparam ii3360.CONFIG_DATA = 16'h5555;
      defparam ii3360.PLACE_LOCATION = "NONE";
      defparam ii3360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3361 ( .DX(nn3361), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2344_), .F2(dummy_abc_2345_), .F3(dummy_abc_2346_) );
      defparam ii3361.CONFIG_DATA = 16'h5555;
      defparam ii3361.PLACE_LOCATION = "NONE";
      defparam ii3361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3362 ( .DX(nn3362), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2347_), .F2(dummy_abc_2348_), .F3(dummy_abc_2349_) );
      defparam ii3362.CONFIG_DATA = 16'h5555;
      defparam ii3362.PLACE_LOCATION = "NONE";
      defparam ii3362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3363 ( .DX(nn3363), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2350_), .F2(dummy_abc_2351_), .F3(dummy_abc_2352_) );
      defparam ii3363.CONFIG_DATA = 16'h5555;
      defparam ii3363.PLACE_LOCATION = "NONE";
      defparam ii3363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3364 ( .DX(nn3364), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2353_), .F2(dummy_abc_2354_), .F3(dummy_abc_2355_) );
      defparam ii3364.CONFIG_DATA = 16'h5555;
      defparam ii3364.PLACE_LOCATION = "NONE";
      defparam ii3364.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_219_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3302, nn3311, nn3309, nn3307, 
              nn3305, nn3347, \coefcal1_xDividend__reg[10]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_151_ ), 
        .DX( {nn3364, nn3363, nn3362, nn3361, nn3360, nn3359, nn3358, nn3357, 
              nn3356, nn3355, nn3354, nn3353, nn3352, nn3351, nn3350, nn3349, 
              nn3348} ), 
        .SUM( {dummy_152_, \coefcal1_divide_inst1_u107_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_14|SUM_net , \coefcal1_divide_inst1_u107_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_12|SUM_net , \coefcal1_divide_inst1_u107_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_10|SUM_net , \coefcal1_divide_inst1_u107_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_8|SUM_net , \coefcal1_divide_inst1_u107_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_6|SUM_net , \coefcal1_divide_inst1_u107_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_4|SUM_net , \coefcal1_divide_inst1_u107_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_2|SUM_net , \coefcal1_divide_inst1_u107_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u107_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3384 ( .DX(nn3384), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_318_), .F2(nn3347), .F3(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ) );
      defparam ii3384.CONFIG_DATA = 16'hA695;
      defparam ii3384.PLACE_LOCATION = "NONE";
      defparam ii3384.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3385 ( .DX(nn3385), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3305), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ) );
      defparam ii3385.CONFIG_DATA = 16'h9A95;
      defparam ii3385.PLACE_LOCATION = "NONE";
      defparam ii3385.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3386 ( .DX(nn3386), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3307), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ) );
      defparam ii3386.CONFIG_DATA = 16'h9A95;
      defparam ii3386.PLACE_LOCATION = "NONE";
      defparam ii3386.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3387 ( .DX(nn3387), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3309), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ) );
      defparam ii3387.CONFIG_DATA = 16'h9A95;
      defparam ii3387.PLACE_LOCATION = "NONE";
      defparam ii3387.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3388 ( .DX(nn3388), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3311), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ) );
      defparam ii3388.CONFIG_DATA = 16'h9A95;
      defparam ii3388.PLACE_LOCATION = "NONE";
      defparam ii3388.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3389 ( .DX(nn3389), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3302), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_6|SUM_net ) );
      defparam ii3389.CONFIG_DATA = 16'h9A95;
      defparam ii3389.PLACE_LOCATION = "NONE";
      defparam ii3389.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3390 ( .DX(nn3390), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2356_), .F2(dummy_abc_2357_), .F3(dummy_abc_2358_) );
      defparam ii3390.CONFIG_DATA = 16'h5555;
      defparam ii3390.PLACE_LOCATION = "NONE";
      defparam ii3390.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3391 ( .DX(nn3391), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2359_), .F2(dummy_abc_2360_), .F3(dummy_abc_2361_) );
      defparam ii3391.CONFIG_DATA = 16'h5555;
      defparam ii3391.PLACE_LOCATION = "NONE";
      defparam ii3391.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3392 ( .DX(nn3392), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2362_), .F2(dummy_abc_2363_), .F3(dummy_abc_2364_) );
      defparam ii3392.CONFIG_DATA = 16'h5555;
      defparam ii3392.PLACE_LOCATION = "NONE";
      defparam ii3392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3393 ( .DX(nn3393), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2365_), .F2(dummy_abc_2366_), .F3(dummy_abc_2367_) );
      defparam ii3393.CONFIG_DATA = 16'h5555;
      defparam ii3393.PLACE_LOCATION = "NONE";
      defparam ii3393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3394 ( .DX(nn3394), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2368_), .F2(dummy_abc_2369_), .F3(dummy_abc_2370_) );
      defparam ii3394.CONFIG_DATA = 16'h5555;
      defparam ii3394.PLACE_LOCATION = "NONE";
      defparam ii3394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3395 ( .DX(nn3395), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2371_), .F2(dummy_abc_2372_), .F3(dummy_abc_2373_) );
      defparam ii3395.CONFIG_DATA = 16'h5555;
      defparam ii3395.PLACE_LOCATION = "NONE";
      defparam ii3395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3396 ( .DX(nn3396), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2374_), .F2(dummy_abc_2375_), .F3(dummy_abc_2376_) );
      defparam ii3396.CONFIG_DATA = 16'h5555;
      defparam ii3396.PLACE_LOCATION = "NONE";
      defparam ii3396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3397 ( .DX(nn3397), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2377_), .F2(dummy_abc_2378_), .F3(dummy_abc_2379_) );
      defparam ii3397.CONFIG_DATA = 16'h5555;
      defparam ii3397.PLACE_LOCATION = "NONE";
      defparam ii3397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3398 ( .DX(nn3398), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2380_), .F2(dummy_abc_2381_), .F3(dummy_abc_2382_) );
      defparam ii3398.CONFIG_DATA = 16'h5555;
      defparam ii3398.PLACE_LOCATION = "NONE";
      defparam ii3398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3399 ( .DX(nn3399), .F0(dummy_abc_2383_), .F1(dummy_abc_2384_), .F2(dummy_abc_2385_), .F3(dummy_abc_2386_) );
      defparam ii3399.CONFIG_DATA = 16'hFFFF;
      defparam ii3399.PLACE_LOCATION = "NONE";
      defparam ii3399.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_235_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_337_ ), 
        .DX( {nn3399, nn3398, nn3397, nn3396, nn3395, nn3394, nn3393, nn3392, 
              nn3391, nn3390, nn3389, nn3388, nn3387, nn3386, nn3385, nn3384, 
              nn3346, nn3345} ), 
        .SUM( {\coefcal1_divide_inst1_u132_XORCI_17|SUM_net , dummy_338_, 
              dummy_339_, dummy_340_, dummy_341_, dummy_342_, dummy_343_, dummy_344_, 
              dummy_345_, dummy_346_, dummy_347_, dummy_348_, dummy_349_, dummy_350_, 
              dummy_351_, dummy_352_, dummy_353_, dummy_354_} )
      );
    CS_LUT4_PRIM ii3420 ( .DX(nn3420), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_318_), .F3(dummy_abc_2387_) );
      defparam ii3420.CONFIG_DATA = 16'hA6A6;
      defparam ii3420.PLACE_LOCATION = "NONE";
      defparam ii3420.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3421 ( .DX(nn3421), .F0(dummy_318_), .F1(nn3347), .F2(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ), .F3(dummy_abc_2388_) );
      defparam ii3421.CONFIG_DATA = 16'hD8D8;
      defparam ii3421.PLACE_LOCATION = "NONE";
      defparam ii3421.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3422 ( .DX(nn3422), .F0(nn3305), .F1(dummy_318_), .F2(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ), .F3(dummy_abc_2389_) );
      defparam ii3422.CONFIG_DATA = 16'hB8B8;
      defparam ii3422.PLACE_LOCATION = "NONE";
      defparam ii3422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3423 ( .DX(nn3423), .F0(nn3307), .F1(dummy_318_), .F2(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ), .F3(dummy_abc_2390_) );
      defparam ii3423.CONFIG_DATA = 16'hB8B8;
      defparam ii3423.PLACE_LOCATION = "NONE";
      defparam ii3423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3424 ( .DX(nn3424), .F0(nn3309), .F1(dummy_318_), .F2(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ), .F3(dummy_abc_2391_) );
      defparam ii3424.CONFIG_DATA = 16'hB8B8;
      defparam ii3424.PLACE_LOCATION = "NONE";
      defparam ii3424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3425 ( .DX(nn3425), .F0(nn3311), .F1(dummy_318_), .F2(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ), .F3(dummy_abc_2392_) );
      defparam ii3425.CONFIG_DATA = 16'hB8B8;
      defparam ii3425.PLACE_LOCATION = "NONE";
      defparam ii3425.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3426 ( .DX(nn3426), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2393_), .F3(dummy_abc_2394_) );
      defparam ii3426.CONFIG_DATA = 16'h9999;
      defparam ii3426.PLACE_LOCATION = "NONE";
      defparam ii3426.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3427 ( .DX(nn3427), .F0(\coefcal1_xDividend__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_318_) );
      defparam ii3427.CONFIG_DATA = 16'hA569;
      defparam ii3427.PLACE_LOCATION = "NONE";
      defparam ii3427.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3428 ( .DX(nn3428), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_318_), .F2(nn3347), .F3(\coefcal1_divide_inst1_u107_XORCI_1|SUM_net ) );
      defparam ii3428.CONFIG_DATA = 16'hA695;
      defparam ii3428.PLACE_LOCATION = "NONE";
      defparam ii3428.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3429 ( .DX(nn3429), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3305), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_2|SUM_net ) );
      defparam ii3429.CONFIG_DATA = 16'h9A95;
      defparam ii3429.PLACE_LOCATION = "NONE";
      defparam ii3429.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3430 ( .DX(nn3430), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3307), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_3|SUM_net ) );
      defparam ii3430.CONFIG_DATA = 16'h9A95;
      defparam ii3430.PLACE_LOCATION = "NONE";
      defparam ii3430.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3431 ( .DX(nn3431), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3309), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_4|SUM_net ) );
      defparam ii3431.CONFIG_DATA = 16'h9A95;
      defparam ii3431.PLACE_LOCATION = "NONE";
      defparam ii3431.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3432 ( .DX(nn3432), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3311), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_5|SUM_net ) );
      defparam ii3432.CONFIG_DATA = 16'h9A95;
      defparam ii3432.PLACE_LOCATION = "NONE";
      defparam ii3432.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3433 ( .DX(nn3433), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3302), .F2(dummy_318_), .F3(\coefcal1_divide_inst1_u107_XORCI_6|SUM_net ) );
      defparam ii3433.CONFIG_DATA = 16'h9A95;
      defparam ii3433.PLACE_LOCATION = "NONE";
      defparam ii3433.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3434 ( .DX(nn3434), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(dummy_abc_2395_), .F2(dummy_abc_2396_), .F3(dummy_abc_2397_) );
      defparam ii3434.CONFIG_DATA = 16'h5555;
      defparam ii3434.PLACE_LOCATION = "NONE";
      defparam ii3434.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3435 ( .DX(nn3435), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2398_), .F2(dummy_abc_2399_), .F3(dummy_abc_2400_) );
      defparam ii3435.CONFIG_DATA = 16'h5555;
      defparam ii3435.PLACE_LOCATION = "NONE";
      defparam ii3435.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3436 ( .DX(nn3436), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2401_), .F2(dummy_abc_2402_), .F3(dummy_abc_2403_) );
      defparam ii3436.CONFIG_DATA = 16'h5555;
      defparam ii3436.PLACE_LOCATION = "NONE";
      defparam ii3436.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3437 ( .DX(nn3437), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2404_), .F2(dummy_abc_2405_), .F3(dummy_abc_2406_) );
      defparam ii3437.CONFIG_DATA = 16'h5555;
      defparam ii3437.PLACE_LOCATION = "NONE";
      defparam ii3437.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3438 ( .DX(nn3438), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2407_), .F2(dummy_abc_2408_), .F3(dummy_abc_2409_) );
      defparam ii3438.CONFIG_DATA = 16'h5555;
      defparam ii3438.PLACE_LOCATION = "NONE";
      defparam ii3438.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3439 ( .DX(nn3439), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2410_), .F2(dummy_abc_2411_), .F3(dummy_abc_2412_) );
      defparam ii3439.CONFIG_DATA = 16'h5555;
      defparam ii3439.PLACE_LOCATION = "NONE";
      defparam ii3439.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3440 ( .DX(nn3440), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2413_), .F2(dummy_abc_2414_), .F3(dummy_abc_2415_) );
      defparam ii3440.CONFIG_DATA = 16'h5555;
      defparam ii3440.PLACE_LOCATION = "NONE";
      defparam ii3440.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3441 ( .DX(nn3441), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2416_), .F2(dummy_abc_2417_), .F3(dummy_abc_2418_) );
      defparam ii3441.CONFIG_DATA = 16'h5555;
      defparam ii3441.PLACE_LOCATION = "NONE";
      defparam ii3441.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3442 ( .DX(nn3442), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2419_), .F2(dummy_abc_2420_), .F3(dummy_abc_2421_) );
      defparam ii3442.CONFIG_DATA = 16'h5555;
      defparam ii3442.PLACE_LOCATION = "NONE";
      defparam ii3442.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_220_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3425, nn3424, nn3423, nn3422, 
              nn3421, nn3420, \coefcal1_xDividend__reg[9]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_153_ ), 
        .DX( {nn3442, nn3441, nn3440, nn3439, nn3438, nn3437, nn3436, nn3435, 
              nn3434, nn3433, nn3432, nn3431, nn3430, nn3429, nn3428, nn3427, 
              nn3426} ), 
        .SUM( {dummy_154_, \coefcal1_divide_inst1_u108_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_14|SUM_net , \coefcal1_divide_inst1_u108_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_12|SUM_net , \coefcal1_divide_inst1_u108_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_10|SUM_net , \coefcal1_divide_inst1_u108_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_8|SUM_net , \coefcal1_divide_inst1_u108_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_6|SUM_net , \coefcal1_divide_inst1_u108_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_4|SUM_net , \coefcal1_divide_inst1_u108_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_2|SUM_net , \coefcal1_divide_inst1_u108_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3462 ( .DX(nn3462), .F0(nn3302), .F1(dummy_318_), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ) );
      defparam ii3462.CONFIG_DATA = 16'h8F80;
      defparam ii3462.PLACE_LOCATION = "NONE";
      defparam ii3462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3463 ( .DX(nn3463), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2422_), .F3(dummy_abc_2423_) );
      defparam ii3463.CONFIG_DATA = 16'h9999;
      defparam ii3463.PLACE_LOCATION = "NONE";
      defparam ii3463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3464 ( .DX(nn3464), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_337_) );
      defparam ii3464.CONFIG_DATA = 16'hA569;
      defparam ii3464.PLACE_LOCATION = "NONE";
      defparam ii3464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3465 ( .DX(nn3465), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_337_), .F2(nn3420), .F3(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ) );
      defparam ii3465.CONFIG_DATA = 16'hA695;
      defparam ii3465.PLACE_LOCATION = "NONE";
      defparam ii3465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3466 ( .DX(nn3466), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3421), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ) );
      defparam ii3466.CONFIG_DATA = 16'h9A95;
      defparam ii3466.PLACE_LOCATION = "NONE";
      defparam ii3466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3467 ( .DX(nn3467), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3422), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ) );
      defparam ii3467.CONFIG_DATA = 16'h9A95;
      defparam ii3467.PLACE_LOCATION = "NONE";
      defparam ii3467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3468 ( .DX(nn3468), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3423), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ) );
      defparam ii3468.CONFIG_DATA = 16'h9A95;
      defparam ii3468.PLACE_LOCATION = "NONE";
      defparam ii3468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3469 ( .DX(nn3469), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3424), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ) );
      defparam ii3469.CONFIG_DATA = 16'h9A95;
      defparam ii3469.PLACE_LOCATION = "NONE";
      defparam ii3469.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3470 ( .DX(nn3470), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3425), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ) );
      defparam ii3470.CONFIG_DATA = 16'h9A95;
      defparam ii3470.PLACE_LOCATION = "NONE";
      defparam ii3470.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3471 ( .DX(nn3471), .F0(nn3302), .F1(dummy_318_), .F2(dummy_abc_2424_), .F3(dummy_abc_2425_) );
      defparam ii3471.CONFIG_DATA = 16'h8888;
      defparam ii3471.PLACE_LOCATION = "NONE";
      defparam ii3471.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3472 ( .DX(nn3472), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3471), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ) );
      defparam ii3472.CONFIG_DATA = 16'h9095;
      defparam ii3472.PLACE_LOCATION = "NONE";
      defparam ii3472.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3473 ( .DX(nn3473), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2426_), .F2(dummy_abc_2427_), .F3(dummy_abc_2428_) );
      defparam ii3473.CONFIG_DATA = 16'h5555;
      defparam ii3473.PLACE_LOCATION = "NONE";
      defparam ii3473.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3474 ( .DX(nn3474), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2429_), .F2(dummy_abc_2430_), .F3(dummy_abc_2431_) );
      defparam ii3474.CONFIG_DATA = 16'h5555;
      defparam ii3474.PLACE_LOCATION = "NONE";
      defparam ii3474.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3475 ( .DX(nn3475), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2432_), .F2(dummy_abc_2433_), .F3(dummy_abc_2434_) );
      defparam ii3475.CONFIG_DATA = 16'h5555;
      defparam ii3475.PLACE_LOCATION = "NONE";
      defparam ii3475.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3476 ( .DX(nn3476), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2435_), .F2(dummy_abc_2436_), .F3(dummy_abc_2437_) );
      defparam ii3476.CONFIG_DATA = 16'h5555;
      defparam ii3476.PLACE_LOCATION = "NONE";
      defparam ii3476.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3477 ( .DX(nn3477), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2438_), .F2(dummy_abc_2439_), .F3(dummy_abc_2440_) );
      defparam ii3477.CONFIG_DATA = 16'h5555;
      defparam ii3477.PLACE_LOCATION = "NONE";
      defparam ii3477.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3478 ( .DX(nn3478), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2441_), .F2(dummy_abc_2442_), .F3(dummy_abc_2443_) );
      defparam ii3478.CONFIG_DATA = 16'h5555;
      defparam ii3478.PLACE_LOCATION = "NONE";
      defparam ii3478.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3479 ( .DX(nn3479), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2444_), .F2(dummy_abc_2445_), .F3(dummy_abc_2446_) );
      defparam ii3479.CONFIG_DATA = 16'h5555;
      defparam ii3479.PLACE_LOCATION = "NONE";
      defparam ii3479.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3480 ( .DX(nn3480), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2447_), .F2(dummy_abc_2448_), .F3(dummy_abc_2449_) );
      defparam ii3480.CONFIG_DATA = 16'h5555;
      defparam ii3480.PLACE_LOCATION = "NONE";
      defparam ii3480.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3481 ( .DX(nn3481), .F0(dummy_abc_2450_), .F1(dummy_abc_2451_), .F2(dummy_abc_2452_), .F3(dummy_abc_2453_) );
      defparam ii3481.CONFIG_DATA = 16'hFFFF;
      defparam ii3481.PLACE_LOCATION = "NONE";
      defparam ii3481.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_236_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_356_ ), 
        .DX( {nn3481, nn3480, nn3479, nn3478, nn3477, nn3476, nn3475, nn3474, 
              nn3473, nn3472, nn3470, nn3469, nn3468, nn3467, nn3466, nn3465, 
              nn3464, nn3463} ), 
        .SUM( {\coefcal1_divide_inst1_u134_XORCI_17|SUM_net , dummy_357_, 
              dummy_358_, dummy_359_, dummy_360_, dummy_361_, dummy_362_, dummy_363_, 
              dummy_364_, dummy_365_, dummy_366_, dummy_367_, dummy_368_, dummy_369_, 
              dummy_370_, dummy_371_, dummy_372_, dummy_373_} )
      );
    CS_LUT4_PRIM ii3502 ( .DX(nn3502), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_337_), .F3(dummy_abc_2454_) );
      defparam ii3502.CONFIG_DATA = 16'hA6A6;
      defparam ii3502.PLACE_LOCATION = "NONE";
      defparam ii3502.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3503 ( .DX(nn3503), .F0(dummy_337_), .F1(nn3420), .F2(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ), .F3(dummy_abc_2455_) );
      defparam ii3503.CONFIG_DATA = 16'hD8D8;
      defparam ii3503.PLACE_LOCATION = "NONE";
      defparam ii3503.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3504 ( .DX(nn3504), .F0(nn3421), .F1(dummy_337_), .F2(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ), .F3(dummy_abc_2456_) );
      defparam ii3504.CONFIG_DATA = 16'hB8B8;
      defparam ii3504.PLACE_LOCATION = "NONE";
      defparam ii3504.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3505 ( .DX(nn3505), .F0(nn3422), .F1(dummy_337_), .F2(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ), .F3(dummy_abc_2457_) );
      defparam ii3505.CONFIG_DATA = 16'hB8B8;
      defparam ii3505.PLACE_LOCATION = "NONE";
      defparam ii3505.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3506 ( .DX(nn3506), .F0(nn3423), .F1(dummy_337_), .F2(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ), .F3(dummy_abc_2458_) );
      defparam ii3506.CONFIG_DATA = 16'hB8B8;
      defparam ii3506.PLACE_LOCATION = "NONE";
      defparam ii3506.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3507 ( .DX(nn3507), .F0(nn3424), .F1(dummy_337_), .F2(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ), .F3(dummy_abc_2459_) );
      defparam ii3507.CONFIG_DATA = 16'hB8B8;
      defparam ii3507.PLACE_LOCATION = "NONE";
      defparam ii3507.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3508 ( .DX(nn3508), .F0(nn3425), .F1(dummy_337_), .F2(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ), .F3(dummy_abc_2460_) );
      defparam ii3508.CONFIG_DATA = 16'hB8B8;
      defparam ii3508.PLACE_LOCATION = "NONE";
      defparam ii3508.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3509 ( .DX(nn3509), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2461_), .F3(dummy_abc_2462_) );
      defparam ii3509.CONFIG_DATA = 16'h9999;
      defparam ii3509.PLACE_LOCATION = "NONE";
      defparam ii3509.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3510 ( .DX(nn3510), .F0(\coefcal1_xDividend__reg[9]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_337_) );
      defparam ii3510.CONFIG_DATA = 16'hA569;
      defparam ii3510.PLACE_LOCATION = "NONE";
      defparam ii3510.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3511 ( .DX(nn3511), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_337_), .F2(nn3420), .F3(\coefcal1_divide_inst1_u108_XORCI_1|SUM_net ) );
      defparam ii3511.CONFIG_DATA = 16'hA695;
      defparam ii3511.PLACE_LOCATION = "NONE";
      defparam ii3511.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3512 ( .DX(nn3512), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3421), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_2|SUM_net ) );
      defparam ii3512.CONFIG_DATA = 16'h9A95;
      defparam ii3512.PLACE_LOCATION = "NONE";
      defparam ii3512.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3513 ( .DX(nn3513), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3422), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_3|SUM_net ) );
      defparam ii3513.CONFIG_DATA = 16'h9A95;
      defparam ii3513.PLACE_LOCATION = "NONE";
      defparam ii3513.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3514 ( .DX(nn3514), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3423), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_4|SUM_net ) );
      defparam ii3514.CONFIG_DATA = 16'h9A95;
      defparam ii3514.PLACE_LOCATION = "NONE";
      defparam ii3514.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3515 ( .DX(nn3515), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3424), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_5|SUM_net ) );
      defparam ii3515.CONFIG_DATA = 16'h9A95;
      defparam ii3515.PLACE_LOCATION = "NONE";
      defparam ii3515.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3516 ( .DX(nn3516), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3425), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_6|SUM_net ) );
      defparam ii3516.CONFIG_DATA = 16'h9A95;
      defparam ii3516.PLACE_LOCATION = "NONE";
      defparam ii3516.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3517 ( .DX(nn3517), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3471), .F2(dummy_337_), .F3(\coefcal1_divide_inst1_u108_XORCI_7|SUM_net ) );
      defparam ii3517.CONFIG_DATA = 16'h9095;
      defparam ii3517.PLACE_LOCATION = "NONE";
      defparam ii3517.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3518 ( .DX(nn3518), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(dummy_abc_2463_), .F2(dummy_abc_2464_), .F3(dummy_abc_2465_) );
      defparam ii3518.CONFIG_DATA = 16'h5555;
      defparam ii3518.PLACE_LOCATION = "NONE";
      defparam ii3518.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3519 ( .DX(nn3519), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2466_), .F2(dummy_abc_2467_), .F3(dummy_abc_2468_) );
      defparam ii3519.CONFIG_DATA = 16'h5555;
      defparam ii3519.PLACE_LOCATION = "NONE";
      defparam ii3519.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3520 ( .DX(nn3520), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2469_), .F2(dummy_abc_2470_), .F3(dummy_abc_2471_) );
      defparam ii3520.CONFIG_DATA = 16'h5555;
      defparam ii3520.PLACE_LOCATION = "NONE";
      defparam ii3520.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3521 ( .DX(nn3521), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2472_), .F2(dummy_abc_2473_), .F3(dummy_abc_2474_) );
      defparam ii3521.CONFIG_DATA = 16'h5555;
      defparam ii3521.PLACE_LOCATION = "NONE";
      defparam ii3521.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3522 ( .DX(nn3522), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2475_), .F2(dummy_abc_2476_), .F3(dummy_abc_2477_) );
      defparam ii3522.CONFIG_DATA = 16'h5555;
      defparam ii3522.PLACE_LOCATION = "NONE";
      defparam ii3522.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3523 ( .DX(nn3523), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2478_), .F2(dummy_abc_2479_), .F3(dummy_abc_2480_) );
      defparam ii3523.CONFIG_DATA = 16'h5555;
      defparam ii3523.PLACE_LOCATION = "NONE";
      defparam ii3523.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3524 ( .DX(nn3524), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2481_), .F2(dummy_abc_2482_), .F3(dummy_abc_2483_) );
      defparam ii3524.CONFIG_DATA = 16'h5555;
      defparam ii3524.PLACE_LOCATION = "NONE";
      defparam ii3524.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3525 ( .DX(nn3525), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2484_), .F2(dummy_abc_2485_), .F3(dummy_abc_2486_) );
      defparam ii3525.CONFIG_DATA = 16'h5555;
      defparam ii3525.PLACE_LOCATION = "NONE";
      defparam ii3525.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_221_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3462, 
              nn3508, nn3507, nn3506, nn3505, nn3504, nn3503, nn3502, 
              \coefcal1_xDividend__reg[8]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_155_ ), 
        .DX( {nn3525, nn3524, nn3523, nn3522, nn3521, nn3520, nn3519, nn3518, 
              nn3517, nn3516, nn3515, nn3514, nn3513, nn3512, nn3511, nn3510, 
              nn3509} ), 
        .SUM( {dummy_156_, \coefcal1_divide_inst1_u109_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_14|SUM_net , \coefcal1_divide_inst1_u109_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_12|SUM_net , \coefcal1_divide_inst1_u109_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_10|SUM_net , \coefcal1_divide_inst1_u109_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_8|SUM_net , \coefcal1_divide_inst1_u109_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_6|SUM_net , \coefcal1_divide_inst1_u109_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_4|SUM_net , \coefcal1_divide_inst1_u109_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_2|SUM_net , \coefcal1_divide_inst1_u109_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u109_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3545 ( .DX(nn3545), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2487_), .F3(dummy_abc_2488_) );
      defparam ii3545.CONFIG_DATA = 16'h9999;
      defparam ii3545.PLACE_LOCATION = "NONE";
      defparam ii3545.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3546 ( .DX(nn3546), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_356_) );
      defparam ii3546.CONFIG_DATA = 16'hA569;
      defparam ii3546.PLACE_LOCATION = "NONE";
      defparam ii3546.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3547 ( .DX(nn3547), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_356_), .F2(nn3502), .F3(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ) );
      defparam ii3547.CONFIG_DATA = 16'hA695;
      defparam ii3547.PLACE_LOCATION = "NONE";
      defparam ii3547.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3548 ( .DX(nn3548), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3503), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ) );
      defparam ii3548.CONFIG_DATA = 16'h9A95;
      defparam ii3548.PLACE_LOCATION = "NONE";
      defparam ii3548.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3549 ( .DX(nn3549), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3504), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ) );
      defparam ii3549.CONFIG_DATA = 16'h9A95;
      defparam ii3549.PLACE_LOCATION = "NONE";
      defparam ii3549.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3550 ( .DX(nn3550), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3505), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ) );
      defparam ii3550.CONFIG_DATA = 16'h9A95;
      defparam ii3550.PLACE_LOCATION = "NONE";
      defparam ii3550.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3551 ( .DX(nn3551), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3506), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ) );
      defparam ii3551.CONFIG_DATA = 16'h9A95;
      defparam ii3551.PLACE_LOCATION = "NONE";
      defparam ii3551.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3552 ( .DX(nn3552), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3507), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ) );
      defparam ii3552.CONFIG_DATA = 16'h9A95;
      defparam ii3552.PLACE_LOCATION = "NONE";
      defparam ii3552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3553 ( .DX(nn3553), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3508), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ) );
      defparam ii3553.CONFIG_DATA = 16'h9A95;
      defparam ii3553.PLACE_LOCATION = "NONE";
      defparam ii3553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3554 ( .DX(nn3554), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3462), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ) );
      defparam ii3554.CONFIG_DATA = 16'h9995;
      defparam ii3554.PLACE_LOCATION = "NONE";
      defparam ii3554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3555 ( .DX(nn3555), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2489_), .F2(dummy_abc_2490_), .F3(dummy_abc_2491_) );
      defparam ii3555.CONFIG_DATA = 16'h5555;
      defparam ii3555.PLACE_LOCATION = "NONE";
      defparam ii3555.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3556 ( .DX(nn3556), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2492_), .F2(dummy_abc_2493_), .F3(dummy_abc_2494_) );
      defparam ii3556.CONFIG_DATA = 16'h5555;
      defparam ii3556.PLACE_LOCATION = "NONE";
      defparam ii3556.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3557 ( .DX(nn3557), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2495_), .F2(dummy_abc_2496_), .F3(dummy_abc_2497_) );
      defparam ii3557.CONFIG_DATA = 16'h5555;
      defparam ii3557.PLACE_LOCATION = "NONE";
      defparam ii3557.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3558 ( .DX(nn3558), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2498_), .F2(dummy_abc_2499_), .F3(dummy_abc_2500_) );
      defparam ii3558.CONFIG_DATA = 16'h5555;
      defparam ii3558.PLACE_LOCATION = "NONE";
      defparam ii3558.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3559 ( .DX(nn3559), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2501_), .F2(dummy_abc_2502_), .F3(dummy_abc_2503_) );
      defparam ii3559.CONFIG_DATA = 16'h5555;
      defparam ii3559.PLACE_LOCATION = "NONE";
      defparam ii3559.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3560 ( .DX(nn3560), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2504_), .F2(dummy_abc_2505_), .F3(dummy_abc_2506_) );
      defparam ii3560.CONFIG_DATA = 16'h5555;
      defparam ii3560.PLACE_LOCATION = "NONE";
      defparam ii3560.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3561 ( .DX(nn3561), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2507_), .F2(dummy_abc_2508_), .F3(dummy_abc_2509_) );
      defparam ii3561.CONFIG_DATA = 16'h5555;
      defparam ii3561.PLACE_LOCATION = "NONE";
      defparam ii3561.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3562 ( .DX(nn3562), .F0(dummy_abc_2510_), .F1(dummy_abc_2511_), .F2(dummy_abc_2512_), .F3(dummy_abc_2513_) );
      defparam ii3562.CONFIG_DATA = 16'hFFFF;
      defparam ii3562.PLACE_LOCATION = "NONE";
      defparam ii3562.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_237_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_375_ ), 
        .DX( {nn3562, nn3561, nn3560, nn3559, nn3558, nn3557, nn3556, nn3555, 
              nn3554, nn3553, nn3552, nn3551, nn3550, nn3549, nn3548, nn3547, 
              nn3546, nn3545} ), 
        .SUM( {\coefcal1_divide_inst1_u136_XORCI_17|SUM_net , dummy_376_, 
              dummy_377_, dummy_378_, dummy_379_, dummy_380_, dummy_381_, dummy_382_, 
              dummy_383_, dummy_384_, dummy_385_, dummy_386_, dummy_387_, dummy_388_, 
              dummy_389_, dummy_390_, dummy_391_, dummy_392_} )
      );
    CS_LUT4_PRIM ii3583 ( .DX(nn3583), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_356_), .F3(dummy_abc_2514_) );
      defparam ii3583.CONFIG_DATA = 16'hA6A6;
      defparam ii3583.PLACE_LOCATION = "NONE";
      defparam ii3583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3584 ( .DX(nn3584), .F0(dummy_356_), .F1(nn3502), .F2(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ), .F3(dummy_abc_2515_) );
      defparam ii3584.CONFIG_DATA = 16'hD8D8;
      defparam ii3584.PLACE_LOCATION = "NONE";
      defparam ii3584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3585 ( .DX(nn3585), .F0(nn3503), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ), .F3(dummy_abc_2516_) );
      defparam ii3585.CONFIG_DATA = 16'hB8B8;
      defparam ii3585.PLACE_LOCATION = "NONE";
      defparam ii3585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3586 ( .DX(nn3586), .F0(nn3504), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ), .F3(dummy_abc_2517_) );
      defparam ii3586.CONFIG_DATA = 16'hB8B8;
      defparam ii3586.PLACE_LOCATION = "NONE";
      defparam ii3586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3587 ( .DX(nn3587), .F0(nn3505), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ), .F3(dummy_abc_2518_) );
      defparam ii3587.CONFIG_DATA = 16'hB8B8;
      defparam ii3587.PLACE_LOCATION = "NONE";
      defparam ii3587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3588 ( .DX(nn3588), .F0(nn3506), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ), .F3(dummy_abc_2519_) );
      defparam ii3588.CONFIG_DATA = 16'hB8B8;
      defparam ii3588.PLACE_LOCATION = "NONE";
      defparam ii3588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3589 ( .DX(nn3589), .F0(nn3507), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ), .F3(dummy_abc_2520_) );
      defparam ii3589.CONFIG_DATA = 16'hB8B8;
      defparam ii3589.PLACE_LOCATION = "NONE";
      defparam ii3589.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3590 ( .DX(nn3590), .F0(nn3508), .F1(dummy_356_), .F2(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ), .F3(dummy_abc_2521_) );
      defparam ii3590.CONFIG_DATA = 16'hB8B8;
      defparam ii3590.PLACE_LOCATION = "NONE";
      defparam ii3590.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3591 ( .DX(nn3591), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2522_), .F3(dummy_abc_2523_) );
      defparam ii3591.CONFIG_DATA = 16'h9999;
      defparam ii3591.PLACE_LOCATION = "NONE";
      defparam ii3591.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3592 ( .DX(nn3592), .F0(\coefcal1_xDividend__reg[8]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_356_) );
      defparam ii3592.CONFIG_DATA = 16'hA569;
      defparam ii3592.PLACE_LOCATION = "NONE";
      defparam ii3592.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3593 ( .DX(nn3593), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_356_), .F2(nn3502), .F3(\coefcal1_divide_inst1_u109_XORCI_1|SUM_net ) );
      defparam ii3593.CONFIG_DATA = 16'hA695;
      defparam ii3593.PLACE_LOCATION = "NONE";
      defparam ii3593.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3594 ( .DX(nn3594), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3503), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_2|SUM_net ) );
      defparam ii3594.CONFIG_DATA = 16'h9A95;
      defparam ii3594.PLACE_LOCATION = "NONE";
      defparam ii3594.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3595 ( .DX(nn3595), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3504), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_3|SUM_net ) );
      defparam ii3595.CONFIG_DATA = 16'h9A95;
      defparam ii3595.PLACE_LOCATION = "NONE";
      defparam ii3595.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3596 ( .DX(nn3596), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3505), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_4|SUM_net ) );
      defparam ii3596.CONFIG_DATA = 16'h9A95;
      defparam ii3596.PLACE_LOCATION = "NONE";
      defparam ii3596.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3597 ( .DX(nn3597), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3506), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_5|SUM_net ) );
      defparam ii3597.CONFIG_DATA = 16'h9A95;
      defparam ii3597.PLACE_LOCATION = "NONE";
      defparam ii3597.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3598 ( .DX(nn3598), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3507), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_6|SUM_net ) );
      defparam ii3598.CONFIG_DATA = 16'h9A95;
      defparam ii3598.PLACE_LOCATION = "NONE";
      defparam ii3598.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3599 ( .DX(nn3599), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3508), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_7|SUM_net ) );
      defparam ii3599.CONFIG_DATA = 16'h9A95;
      defparam ii3599.PLACE_LOCATION = "NONE";
      defparam ii3599.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3600 ( .DX(nn3600), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3462), .F2(dummy_356_), .F3(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ) );
      defparam ii3600.CONFIG_DATA = 16'h9995;
      defparam ii3600.PLACE_LOCATION = "NONE";
      defparam ii3600.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3601 ( .DX(nn3601), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(dummy_abc_2524_), .F2(dummy_abc_2525_), .F3(dummy_abc_2526_) );
      defparam ii3601.CONFIG_DATA = 16'h5555;
      defparam ii3601.PLACE_LOCATION = "NONE";
      defparam ii3601.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3602 ( .DX(nn3602), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2527_), .F2(dummy_abc_2528_), .F3(dummy_abc_2529_) );
      defparam ii3602.CONFIG_DATA = 16'h5555;
      defparam ii3602.PLACE_LOCATION = "NONE";
      defparam ii3602.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3603 ( .DX(nn3603), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2530_), .F2(dummy_abc_2531_), .F3(dummy_abc_2532_) );
      defparam ii3603.CONFIG_DATA = 16'h5555;
      defparam ii3603.PLACE_LOCATION = "NONE";
      defparam ii3603.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3604 ( .DX(nn3604), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2533_), .F2(dummy_abc_2534_), .F3(dummy_abc_2535_) );
      defparam ii3604.CONFIG_DATA = 16'h5555;
      defparam ii3604.PLACE_LOCATION = "NONE";
      defparam ii3604.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3605 ( .DX(nn3605), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2536_), .F2(dummy_abc_2537_), .F3(dummy_abc_2538_) );
      defparam ii3605.CONFIG_DATA = 16'h5555;
      defparam ii3605.PLACE_LOCATION = "NONE";
      defparam ii3605.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3606 ( .DX(nn3606), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2539_), .F2(dummy_abc_2540_), .F3(dummy_abc_2541_) );
      defparam ii3606.CONFIG_DATA = 16'h5555;
      defparam ii3606.PLACE_LOCATION = "NONE";
      defparam ii3606.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3607 ( .DX(nn3607), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2542_), .F2(dummy_abc_2543_), .F3(dummy_abc_2544_) );
      defparam ii3607.CONFIG_DATA = 16'h5555;
      defparam ii3607.PLACE_LOCATION = "NONE";
      defparam ii3607.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_222_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3590, 
              nn3589, nn3588, nn3587, nn3586, nn3585, nn3584, nn3583, 
              \coefcal1_xDividend__reg[7]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_157_ ), 
        .DX( {nn3607, nn3606, nn3605, nn3604, nn3603, nn3602, nn3601, nn3600, 
              nn3599, nn3598, nn3597, nn3596, nn3595, nn3594, nn3593, nn3592, 
              nn3591} ), 
        .SUM( {dummy_158_, \coefcal1_divide_inst1_u110_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_14|SUM_net , \coefcal1_divide_inst1_u110_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_12|SUM_net , \coefcal1_divide_inst1_u110_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_10|SUM_net , \coefcal1_divide_inst1_u110_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_8|SUM_net , \coefcal1_divide_inst1_u110_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_6|SUM_net , \coefcal1_divide_inst1_u110_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_4|SUM_net , \coefcal1_divide_inst1_u110_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_2|SUM_net , \coefcal1_divide_inst1_u110_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3627 ( .DX(nn3627), .F0(dummy_356_), .F1(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ), .F2(dummy_375_), .F3(\coefcal1_divide_inst1_u110_XORCI_9|SUM_net ) );
      defparam ii3627.CONFIG_DATA = 16'hEFE0;
      defparam ii3627.PLACE_LOCATION = "NONE";
      defparam ii3627.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3628 ( .DX(nn3628), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2545_), .F3(dummy_abc_2546_) );
      defparam ii3628.CONFIG_DATA = 16'h9999;
      defparam ii3628.PLACE_LOCATION = "NONE";
      defparam ii3628.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3629 ( .DX(nn3629), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_375_) );
      defparam ii3629.CONFIG_DATA = 16'hA569;
      defparam ii3629.PLACE_LOCATION = "NONE";
      defparam ii3629.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3630 ( .DX(nn3630), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_375_), .F2(nn3583), .F3(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ) );
      defparam ii3630.CONFIG_DATA = 16'hA695;
      defparam ii3630.PLACE_LOCATION = "NONE";
      defparam ii3630.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3631 ( .DX(nn3631), .F0(nn3584), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_2|SUM_net ), .F3(dummy_abc_2547_) );
      defparam ii3631.CONFIG_DATA = 16'hB8B8;
      defparam ii3631.PLACE_LOCATION = "NONE";
      defparam ii3631.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3632 ( .DX(nn3632), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3631), .F2(dummy_abc_2548_), .F3(dummy_abc_2549_) );
      defparam ii3632.CONFIG_DATA = 16'h9999;
      defparam ii3632.PLACE_LOCATION = "NONE";
      defparam ii3632.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3633 ( .DX(nn3633), .F0(nn3585), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_3|SUM_net ), .F3(dummy_abc_2550_) );
      defparam ii3633.CONFIG_DATA = 16'hB8B8;
      defparam ii3633.PLACE_LOCATION = "NONE";
      defparam ii3633.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3634 ( .DX(nn3634), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3633), .F2(dummy_abc_2551_), .F3(dummy_abc_2552_) );
      defparam ii3634.CONFIG_DATA = 16'h9999;
      defparam ii3634.PLACE_LOCATION = "NONE";
      defparam ii3634.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3635 ( .DX(nn3635), .F0(nn3586), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_4|SUM_net ), .F3(dummy_abc_2553_) );
      defparam ii3635.CONFIG_DATA = 16'hB8B8;
      defparam ii3635.PLACE_LOCATION = "NONE";
      defparam ii3635.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3636 ( .DX(nn3636), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3635), .F2(dummy_abc_2554_), .F3(dummy_abc_2555_) );
      defparam ii3636.CONFIG_DATA = 16'h9999;
      defparam ii3636.PLACE_LOCATION = "NONE";
      defparam ii3636.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3637 ( .DX(nn3637), .F0(nn3587), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_5|SUM_net ), .F3(dummy_abc_2556_) );
      defparam ii3637.CONFIG_DATA = 16'hB8B8;
      defparam ii3637.PLACE_LOCATION = "NONE";
      defparam ii3637.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3638 ( .DX(nn3638), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3637), .F2(dummy_abc_2557_), .F3(dummy_abc_2558_) );
      defparam ii3638.CONFIG_DATA = 16'h9999;
      defparam ii3638.PLACE_LOCATION = "NONE";
      defparam ii3638.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3639 ( .DX(nn3639), .F0(nn3588), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_6|SUM_net ), .F3(dummy_abc_2559_) );
      defparam ii3639.CONFIG_DATA = 16'hB8B8;
      defparam ii3639.PLACE_LOCATION = "NONE";
      defparam ii3639.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3640 ( .DX(nn3640), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3639), .F2(dummy_abc_2560_), .F3(dummy_abc_2561_) );
      defparam ii3640.CONFIG_DATA = 16'h9999;
      defparam ii3640.PLACE_LOCATION = "NONE";
      defparam ii3640.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3641 ( .DX(nn3641), .F0(nn3589), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_7|SUM_net ), .F3(dummy_abc_2562_) );
      defparam ii3641.CONFIG_DATA = 16'hB8B8;
      defparam ii3641.PLACE_LOCATION = "NONE";
      defparam ii3641.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3642 ( .DX(nn3642), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3641), .F2(dummy_abc_2563_), .F3(dummy_abc_2564_) );
      defparam ii3642.CONFIG_DATA = 16'h9999;
      defparam ii3642.PLACE_LOCATION = "NONE";
      defparam ii3642.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3643 ( .DX(nn3643), .F0(nn3590), .F1(dummy_375_), .F2(\coefcal1_divide_inst1_u110_XORCI_8|SUM_net ), .F3(dummy_abc_2565_) );
      defparam ii3643.CONFIG_DATA = 16'hB8B8;
      defparam ii3643.PLACE_LOCATION = "NONE";
      defparam ii3643.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3644 ( .DX(nn3644), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3643), .F2(dummy_abc_2566_), .F3(dummy_abc_2567_) );
      defparam ii3644.CONFIG_DATA = 16'h9999;
      defparam ii3644.PLACE_LOCATION = "NONE";
      defparam ii3644.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3645 ( .DX(nn3645), .F0(dummy_356_), .F1(\coefcal1_divide_inst1_u109_XORCI_8|SUM_net ), .F2(dummy_abc_2568_), .F3(dummy_abc_2569_) );
      defparam ii3645.CONFIG_DATA = 16'h1111;
      defparam ii3645.PLACE_LOCATION = "NONE";
      defparam ii3645.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3646 ( .DX(nn3646), .F0(nn3462), .F1(nn3645), .F2(dummy_375_), .F3(\coefcal1_divide_inst1_u110_XORCI_9|SUM_net ) );
      defparam ii3646.CONFIG_DATA = 16'h2A20;
      defparam ii3646.PLACE_LOCATION = "NONE";
      defparam ii3646.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3647 ( .DX(nn3647), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3646), .F2(dummy_abc_2570_), .F3(dummy_abc_2571_) );
      defparam ii3647.CONFIG_DATA = 16'h9999;
      defparam ii3647.PLACE_LOCATION = "NONE";
      defparam ii3647.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3648 ( .DX(nn3648), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2572_), .F2(dummy_abc_2573_), .F3(dummy_abc_2574_) );
      defparam ii3648.CONFIG_DATA = 16'h5555;
      defparam ii3648.PLACE_LOCATION = "NONE";
      defparam ii3648.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3649 ( .DX(nn3649), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2575_), .F2(dummy_abc_2576_), .F3(dummy_abc_2577_) );
      defparam ii3649.CONFIG_DATA = 16'h5555;
      defparam ii3649.PLACE_LOCATION = "NONE";
      defparam ii3649.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3650 ( .DX(nn3650), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2578_), .F2(dummy_abc_2579_), .F3(dummy_abc_2580_) );
      defparam ii3650.CONFIG_DATA = 16'h5555;
      defparam ii3650.PLACE_LOCATION = "NONE";
      defparam ii3650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3651 ( .DX(nn3651), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2581_), .F2(dummy_abc_2582_), .F3(dummy_abc_2583_) );
      defparam ii3651.CONFIG_DATA = 16'h5555;
      defparam ii3651.PLACE_LOCATION = "NONE";
      defparam ii3651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3652 ( .DX(nn3652), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2584_), .F2(dummy_abc_2585_), .F3(dummy_abc_2586_) );
      defparam ii3652.CONFIG_DATA = 16'h5555;
      defparam ii3652.PLACE_LOCATION = "NONE";
      defparam ii3652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3653 ( .DX(nn3653), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2587_), .F2(dummy_abc_2588_), .F3(dummy_abc_2589_) );
      defparam ii3653.CONFIG_DATA = 16'h5555;
      defparam ii3653.PLACE_LOCATION = "NONE";
      defparam ii3653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3654 ( .DX(nn3654), .F0(dummy_abc_2590_), .F1(dummy_abc_2591_), .F2(dummy_abc_2592_), .F3(dummy_abc_2593_) );
      defparam ii3654.CONFIG_DATA = 16'hFFFF;
      defparam ii3654.PLACE_LOCATION = "NONE";
      defparam ii3654.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_238_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_394_ ), 
        .DX( {nn3654, nn3653, nn3652, nn3651, nn3650, nn3649, nn3648, nn3647, 
              nn3644, nn3642, nn3640, nn3638, nn3636, nn3634, nn3632, nn3630, 
              nn3629, nn3628} ), 
        .SUM( {\coefcal1_divide_inst1_u138_XORCI_17|SUM_net , dummy_395_, 
              dummy_396_, dummy_397_, dummy_398_, dummy_399_, dummy_400_, dummy_401_, 
              dummy_402_, dummy_403_, dummy_404_, dummy_405_, dummy_406_, dummy_407_, 
              dummy_408_, dummy_409_, dummy_410_, dummy_411_} )
      );
    CS_LUT4_PRIM ii3675 ( .DX(nn3675), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_375_), .F3(dummy_abc_2594_) );
      defparam ii3675.CONFIG_DATA = 16'hA6A6;
      defparam ii3675.PLACE_LOCATION = "NONE";
      defparam ii3675.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3676 ( .DX(nn3676), .F0(dummy_375_), .F1(nn3583), .F2(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ), .F3(dummy_abc_2595_) );
      defparam ii3676.CONFIG_DATA = 16'hD8D8;
      defparam ii3676.PLACE_LOCATION = "NONE";
      defparam ii3676.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3677 ( .DX(nn3677), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2596_), .F3(dummy_abc_2597_) );
      defparam ii3677.CONFIG_DATA = 16'h9999;
      defparam ii3677.PLACE_LOCATION = "NONE";
      defparam ii3677.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3678 ( .DX(nn3678), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_375_) );
      defparam ii3678.CONFIG_DATA = 16'hA569;
      defparam ii3678.PLACE_LOCATION = "NONE";
      defparam ii3678.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3679 ( .DX(nn3679), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_375_), .F2(nn3583), .F3(\coefcal1_divide_inst1_u110_XORCI_1|SUM_net ) );
      defparam ii3679.CONFIG_DATA = 16'hA695;
      defparam ii3679.PLACE_LOCATION = "NONE";
      defparam ii3679.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3680 ( .DX(nn3680), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3631), .F2(dummy_abc_2598_), .F3(dummy_abc_2599_) );
      defparam ii3680.CONFIG_DATA = 16'h9999;
      defparam ii3680.PLACE_LOCATION = "NONE";
      defparam ii3680.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3681 ( .DX(nn3681), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3633), .F2(dummy_abc_2600_), .F3(dummy_abc_2601_) );
      defparam ii3681.CONFIG_DATA = 16'h9999;
      defparam ii3681.PLACE_LOCATION = "NONE";
      defparam ii3681.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3682 ( .DX(nn3682), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3635), .F2(dummy_abc_2602_), .F3(dummy_abc_2603_) );
      defparam ii3682.CONFIG_DATA = 16'h9999;
      defparam ii3682.PLACE_LOCATION = "NONE";
      defparam ii3682.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3683 ( .DX(nn3683), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3637), .F2(dummy_abc_2604_), .F3(dummy_abc_2605_) );
      defparam ii3683.CONFIG_DATA = 16'h9999;
      defparam ii3683.PLACE_LOCATION = "NONE";
      defparam ii3683.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3684 ( .DX(nn3684), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3639), .F2(dummy_abc_2606_), .F3(dummy_abc_2607_) );
      defparam ii3684.CONFIG_DATA = 16'h9999;
      defparam ii3684.PLACE_LOCATION = "NONE";
      defparam ii3684.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3685 ( .DX(nn3685), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3641), .F2(dummy_abc_2608_), .F3(dummy_abc_2609_) );
      defparam ii3685.CONFIG_DATA = 16'h9999;
      defparam ii3685.PLACE_LOCATION = "NONE";
      defparam ii3685.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3686 ( .DX(nn3686), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3643), .F2(dummy_abc_2610_), .F3(dummy_abc_2611_) );
      defparam ii3686.CONFIG_DATA = 16'h9999;
      defparam ii3686.PLACE_LOCATION = "NONE";
      defparam ii3686.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3687 ( .DX(nn3687), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3646), .F2(dummy_abc_2612_), .F3(dummy_abc_2613_) );
      defparam ii3687.CONFIG_DATA = 16'h9999;
      defparam ii3687.PLACE_LOCATION = "NONE";
      defparam ii3687.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3688 ( .DX(nn3688), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(dummy_abc_2614_), .F2(dummy_abc_2615_), .F3(dummy_abc_2616_) );
      defparam ii3688.CONFIG_DATA = 16'h5555;
      defparam ii3688.PLACE_LOCATION = "NONE";
      defparam ii3688.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3689 ( .DX(nn3689), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2617_), .F2(dummy_abc_2618_), .F3(dummy_abc_2619_) );
      defparam ii3689.CONFIG_DATA = 16'h5555;
      defparam ii3689.PLACE_LOCATION = "NONE";
      defparam ii3689.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3690 ( .DX(nn3690), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2620_), .F2(dummy_abc_2621_), .F3(dummy_abc_2622_) );
      defparam ii3690.CONFIG_DATA = 16'h5555;
      defparam ii3690.PLACE_LOCATION = "NONE";
      defparam ii3690.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3691 ( .DX(nn3691), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2623_), .F2(dummy_abc_2624_), .F3(dummy_abc_2625_) );
      defparam ii3691.CONFIG_DATA = 16'h5555;
      defparam ii3691.PLACE_LOCATION = "NONE";
      defparam ii3691.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3692 ( .DX(nn3692), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2626_), .F2(dummy_abc_2627_), .F3(dummy_abc_2628_) );
      defparam ii3692.CONFIG_DATA = 16'h5555;
      defparam ii3692.PLACE_LOCATION = "NONE";
      defparam ii3692.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3693 ( .DX(nn3693), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2629_), .F2(dummy_abc_2630_), .F3(dummy_abc_2631_) );
      defparam ii3693.CONFIG_DATA = 16'h5555;
      defparam ii3693.PLACE_LOCATION = "NONE";
      defparam ii3693.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_223_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn3646, nn3643, nn3641, nn3639, nn3637, nn3635, nn3633, 
              nn3631, nn3676, nn3675, \coefcal1_xDividend__reg[6]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_159_ ), 
        .DX( {nn3693, nn3692, nn3691, nn3690, nn3689, nn3688, nn3687, nn3686, 
              nn3685, nn3684, nn3683, nn3682, nn3681, nn3680, nn3679, nn3678, 
              nn3677} ), 
        .SUM( {dummy_160_, \coefcal1_divide_inst1_u111_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_14|SUM_net , \coefcal1_divide_inst1_u111_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_12|SUM_net , \coefcal1_divide_inst1_u111_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_10|SUM_net , \coefcal1_divide_inst1_u111_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_8|SUM_net , \coefcal1_divide_inst1_u111_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_6|SUM_net , \coefcal1_divide_inst1_u111_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_4|SUM_net , \coefcal1_divide_inst1_u111_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_2|SUM_net , \coefcal1_divide_inst1_u111_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3713 ( .DX(nn3713), .F0(nn3462), .F1(nn3627), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_10|SUM_net ) );
      defparam ii3713.CONFIG_DATA = 16'h8A80;
      defparam ii3713.PLACE_LOCATION = "NONE";
      defparam ii3713.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3714 ( .DX(nn3714), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2632_), .F3(dummy_abc_2633_) );
      defparam ii3714.CONFIG_DATA = 16'h9999;
      defparam ii3714.PLACE_LOCATION = "NONE";
      defparam ii3714.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3715 ( .DX(nn3715), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_394_) );
      defparam ii3715.CONFIG_DATA = 16'hA569;
      defparam ii3715.PLACE_LOCATION = "NONE";
      defparam ii3715.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3716 ( .DX(nn3716), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_394_), .F2(nn3675), .F3(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ) );
      defparam ii3716.CONFIG_DATA = 16'hA695;
      defparam ii3716.PLACE_LOCATION = "NONE";
      defparam ii3716.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3717 ( .DX(nn3717), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3676), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ) );
      defparam ii3717.CONFIG_DATA = 16'h9A95;
      defparam ii3717.PLACE_LOCATION = "NONE";
      defparam ii3717.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3718 ( .DX(nn3718), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3631), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ) );
      defparam ii3718.CONFIG_DATA = 16'h9A95;
      defparam ii3718.PLACE_LOCATION = "NONE";
      defparam ii3718.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3719 ( .DX(nn3719), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3633), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ) );
      defparam ii3719.CONFIG_DATA = 16'h9A95;
      defparam ii3719.PLACE_LOCATION = "NONE";
      defparam ii3719.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3720 ( .DX(nn3720), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3635), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ) );
      defparam ii3720.CONFIG_DATA = 16'h9A95;
      defparam ii3720.PLACE_LOCATION = "NONE";
      defparam ii3720.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3721 ( .DX(nn3721), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3637), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ) );
      defparam ii3721.CONFIG_DATA = 16'h9A95;
      defparam ii3721.PLACE_LOCATION = "NONE";
      defparam ii3721.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3722 ( .DX(nn3722), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3639), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ) );
      defparam ii3722.CONFIG_DATA = 16'h9A95;
      defparam ii3722.PLACE_LOCATION = "NONE";
      defparam ii3722.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3723 ( .DX(nn3723), .F0(nn3641), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_8|SUM_net ), .F3(dummy_abc_2634_) );
      defparam ii3723.CONFIG_DATA = 16'hB8B8;
      defparam ii3723.PLACE_LOCATION = "NONE";
      defparam ii3723.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3724 ( .DX(nn3724), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3723), .F2(dummy_abc_2635_), .F3(dummy_abc_2636_) );
      defparam ii3724.CONFIG_DATA = 16'h9999;
      defparam ii3724.PLACE_LOCATION = "NONE";
      defparam ii3724.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3725 ( .DX(nn3725), .F0(nn3643), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_9|SUM_net ), .F3(dummy_abc_2637_) );
      defparam ii3725.CONFIG_DATA = 16'hB8B8;
      defparam ii3725.PLACE_LOCATION = "NONE";
      defparam ii3725.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3726 ( .DX(nn3726), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3725), .F2(dummy_abc_2638_), .F3(dummy_abc_2639_) );
      defparam ii3726.CONFIG_DATA = 16'h9999;
      defparam ii3726.PLACE_LOCATION = "NONE";
      defparam ii3726.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3727 ( .DX(nn3727), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3713), .F2(dummy_abc_2640_), .F3(dummy_abc_2641_) );
      defparam ii3727.CONFIG_DATA = 16'h9999;
      defparam ii3727.PLACE_LOCATION = "NONE";
      defparam ii3727.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3728 ( .DX(nn3728), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2642_), .F2(dummy_abc_2643_), .F3(dummy_abc_2644_) );
      defparam ii3728.CONFIG_DATA = 16'h5555;
      defparam ii3728.PLACE_LOCATION = "NONE";
      defparam ii3728.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3729 ( .DX(nn3729), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2645_), .F2(dummy_abc_2646_), .F3(dummy_abc_2647_) );
      defparam ii3729.CONFIG_DATA = 16'h5555;
      defparam ii3729.PLACE_LOCATION = "NONE";
      defparam ii3729.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3730 ( .DX(nn3730), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2648_), .F2(dummy_abc_2649_), .F3(dummy_abc_2650_) );
      defparam ii3730.CONFIG_DATA = 16'h5555;
      defparam ii3730.PLACE_LOCATION = "NONE";
      defparam ii3730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3731 ( .DX(nn3731), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2651_), .F2(dummy_abc_2652_), .F3(dummy_abc_2653_) );
      defparam ii3731.CONFIG_DATA = 16'h5555;
      defparam ii3731.PLACE_LOCATION = "NONE";
      defparam ii3731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3732 ( .DX(nn3732), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2654_), .F2(dummy_abc_2655_), .F3(dummy_abc_2656_) );
      defparam ii3732.CONFIG_DATA = 16'h5555;
      defparam ii3732.PLACE_LOCATION = "NONE";
      defparam ii3732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3733 ( .DX(nn3733), .F0(dummy_abc_2657_), .F1(dummy_abc_2658_), .F2(dummy_abc_2659_), .F3(dummy_abc_2660_) );
      defparam ii3733.CONFIG_DATA = 16'hFFFF;
      defparam ii3733.PLACE_LOCATION = "NONE";
      defparam ii3733.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_239_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_413_ ), 
        .DX( {nn3733, nn3732, nn3731, nn3730, nn3729, nn3728, nn3727, nn3726, 
              nn3724, nn3722, nn3721, nn3720, nn3719, nn3718, nn3717, nn3716, 
              nn3715, nn3714} ), 
        .SUM( {\coefcal1_divide_inst1_u140_XORCI_17|SUM_net , dummy_414_, 
              dummy_415_, dummy_416_, dummy_417_, dummy_418_, dummy_419_, dummy_420_, 
              dummy_421_, dummy_422_, dummy_423_, dummy_424_, dummy_425_, dummy_426_, 
              dummy_427_, dummy_428_, dummy_429_, dummy_430_} )
      );
    CS_LUT4_PRIM ii3754 ( .DX(nn3754), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2661_), .F3(dummy_abc_2662_) );
      defparam ii3754.CONFIG_DATA = 16'h9999;
      defparam ii3754.PLACE_LOCATION = "NONE";
      defparam ii3754.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3755 ( .DX(nn3755), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_413_) );
      defparam ii3755.CONFIG_DATA = 16'hA569;
      defparam ii3755.PLACE_LOCATION = "NONE";
      defparam ii3755.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3756 ( .DX(nn3756), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_394_), .F3(dummy_abc_2663_) );
      defparam ii3756.CONFIG_DATA = 16'hA6A6;
      defparam ii3756.PLACE_LOCATION = "NONE";
      defparam ii3756.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3757 ( .DX(nn3757), .F0(dummy_394_), .F1(nn3675), .F2(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ), .F3(dummy_abc_2664_) );
      defparam ii3757.CONFIG_DATA = 16'hD8D8;
      defparam ii3757.PLACE_LOCATION = "NONE";
      defparam ii3757.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3758 ( .DX(nn3758), .F0(nn3676), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ), .F3(dummy_abc_2665_) );
      defparam ii3758.CONFIG_DATA = 16'hB8B8;
      defparam ii3758.PLACE_LOCATION = "NONE";
      defparam ii3758.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3759 ( .DX(nn3759), .F0(nn3631), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ), .F3(dummy_abc_2666_) );
      defparam ii3759.CONFIG_DATA = 16'hB8B8;
      defparam ii3759.PLACE_LOCATION = "NONE";
      defparam ii3759.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3760 ( .DX(nn3760), .F0(nn3633), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ), .F3(dummy_abc_2667_) );
      defparam ii3760.CONFIG_DATA = 16'hB8B8;
      defparam ii3760.PLACE_LOCATION = "NONE";
      defparam ii3760.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3761 ( .DX(nn3761), .F0(nn3635), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ), .F3(dummy_abc_2668_) );
      defparam ii3761.CONFIG_DATA = 16'hB8B8;
      defparam ii3761.PLACE_LOCATION = "NONE";
      defparam ii3761.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3762 ( .DX(nn3762), .F0(nn3637), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ), .F3(dummy_abc_2669_) );
      defparam ii3762.CONFIG_DATA = 16'hB8B8;
      defparam ii3762.PLACE_LOCATION = "NONE";
      defparam ii3762.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3763 ( .DX(nn3763), .F0(nn3639), .F1(dummy_394_), .F2(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ), .F3(dummy_abc_2670_) );
      defparam ii3763.CONFIG_DATA = 16'hB8B8;
      defparam ii3763.PLACE_LOCATION = "NONE";
      defparam ii3763.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3764 ( .DX(nn3764), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2671_), .F3(dummy_abc_2672_) );
      defparam ii3764.CONFIG_DATA = 16'h9999;
      defparam ii3764.PLACE_LOCATION = "NONE";
      defparam ii3764.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3765 ( .DX(nn3765), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_394_) );
      defparam ii3765.CONFIG_DATA = 16'hA569;
      defparam ii3765.PLACE_LOCATION = "NONE";
      defparam ii3765.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3766 ( .DX(nn3766), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_394_), .F2(nn3675), .F3(\coefcal1_divide_inst1_u111_XORCI_1|SUM_net ) );
      defparam ii3766.CONFIG_DATA = 16'hA695;
      defparam ii3766.PLACE_LOCATION = "NONE";
      defparam ii3766.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3767 ( .DX(nn3767), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3676), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_2|SUM_net ) );
      defparam ii3767.CONFIG_DATA = 16'h9A95;
      defparam ii3767.PLACE_LOCATION = "NONE";
      defparam ii3767.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3768 ( .DX(nn3768), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3631), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_3|SUM_net ) );
      defparam ii3768.CONFIG_DATA = 16'h9A95;
      defparam ii3768.PLACE_LOCATION = "NONE";
      defparam ii3768.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3769 ( .DX(nn3769), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3633), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_4|SUM_net ) );
      defparam ii3769.CONFIG_DATA = 16'h9A95;
      defparam ii3769.PLACE_LOCATION = "NONE";
      defparam ii3769.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3770 ( .DX(nn3770), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3635), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_5|SUM_net ) );
      defparam ii3770.CONFIG_DATA = 16'h9A95;
      defparam ii3770.PLACE_LOCATION = "NONE";
      defparam ii3770.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3771 ( .DX(nn3771), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3637), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_6|SUM_net ) );
      defparam ii3771.CONFIG_DATA = 16'h9A95;
      defparam ii3771.PLACE_LOCATION = "NONE";
      defparam ii3771.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3772 ( .DX(nn3772), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3639), .F2(dummy_394_), .F3(\coefcal1_divide_inst1_u111_XORCI_7|SUM_net ) );
      defparam ii3772.CONFIG_DATA = 16'h9A95;
      defparam ii3772.PLACE_LOCATION = "NONE";
      defparam ii3772.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3773 ( .DX(nn3773), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3723), .F2(dummy_abc_2673_), .F3(dummy_abc_2674_) );
      defparam ii3773.CONFIG_DATA = 16'h9999;
      defparam ii3773.PLACE_LOCATION = "NONE";
      defparam ii3773.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3774 ( .DX(nn3774), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3725), .F2(dummy_abc_2675_), .F3(dummy_abc_2676_) );
      defparam ii3774.CONFIG_DATA = 16'h9999;
      defparam ii3774.PLACE_LOCATION = "NONE";
      defparam ii3774.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3775 ( .DX(nn3775), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3713), .F2(dummy_abc_2677_), .F3(dummy_abc_2678_) );
      defparam ii3775.CONFIG_DATA = 16'h9999;
      defparam ii3775.PLACE_LOCATION = "NONE";
      defparam ii3775.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3776 ( .DX(nn3776), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(dummy_abc_2679_), .F2(dummy_abc_2680_), .F3(dummy_abc_2681_) );
      defparam ii3776.CONFIG_DATA = 16'h5555;
      defparam ii3776.PLACE_LOCATION = "NONE";
      defparam ii3776.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3777 ( .DX(nn3777), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2682_), .F2(dummy_abc_2683_), .F3(dummy_abc_2684_) );
      defparam ii3777.CONFIG_DATA = 16'h5555;
      defparam ii3777.PLACE_LOCATION = "NONE";
      defparam ii3777.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3778 ( .DX(nn3778), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2685_), .F2(dummy_abc_2686_), .F3(dummy_abc_2687_) );
      defparam ii3778.CONFIG_DATA = 16'h5555;
      defparam ii3778.PLACE_LOCATION = "NONE";
      defparam ii3778.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3779 ( .DX(nn3779), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2688_), .F2(dummy_abc_2689_), .F3(dummy_abc_2690_) );
      defparam ii3779.CONFIG_DATA = 16'h5555;
      defparam ii3779.PLACE_LOCATION = "NONE";
      defparam ii3779.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3780 ( .DX(nn3780), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2691_), .F2(dummy_abc_2692_), .F3(dummy_abc_2693_) );
      defparam ii3780.CONFIG_DATA = 16'h5555;
      defparam ii3780.PLACE_LOCATION = "NONE";
      defparam ii3780.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_224_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3713, 
              nn3725, nn3723, nn3763, nn3762, nn3761, nn3760, nn3759, nn3758, 
              nn3757, nn3756, \coefcal1_xDividend__reg[5]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_161_ ), 
        .DX( {nn3780, nn3779, nn3778, nn3777, nn3776, nn3775, nn3774, nn3773, 
              nn3772, nn3771, nn3770, nn3769, nn3768, nn3767, nn3766, nn3765, 
              nn3764} ), 
        .SUM( {dummy_162_, \coefcal1_divide_inst1_u112_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_14|SUM_net , \coefcal1_divide_inst1_u112_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_12|SUM_net , \coefcal1_divide_inst1_u112_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_10|SUM_net , \coefcal1_divide_inst1_u112_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_8|SUM_net , \coefcal1_divide_inst1_u112_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_6|SUM_net , \coefcal1_divide_inst1_u112_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_4|SUM_net , \coefcal1_divide_inst1_u112_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_2|SUM_net , \coefcal1_divide_inst1_u112_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3800 ( .DX(nn3800), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_413_), .F2(nn3756), .F3(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ) );
      defparam ii3800.CONFIG_DATA = 16'hA695;
      defparam ii3800.PLACE_LOCATION = "NONE";
      defparam ii3800.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3801 ( .DX(nn3801), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3757), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ) );
      defparam ii3801.CONFIG_DATA = 16'h9A95;
      defparam ii3801.PLACE_LOCATION = "NONE";
      defparam ii3801.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3802 ( .DX(nn3802), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3758), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ) );
      defparam ii3802.CONFIG_DATA = 16'h9A95;
      defparam ii3802.PLACE_LOCATION = "NONE";
      defparam ii3802.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3803 ( .DX(nn3803), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3759), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ) );
      defparam ii3803.CONFIG_DATA = 16'h9A95;
      defparam ii3803.PLACE_LOCATION = "NONE";
      defparam ii3803.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3804 ( .DX(nn3804), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3760), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ) );
      defparam ii3804.CONFIG_DATA = 16'h9A95;
      defparam ii3804.PLACE_LOCATION = "NONE";
      defparam ii3804.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3805 ( .DX(nn3805), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3761), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ) );
      defparam ii3805.CONFIG_DATA = 16'h9A95;
      defparam ii3805.PLACE_LOCATION = "NONE";
      defparam ii3805.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3806 ( .DX(nn3806), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3762), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ) );
      defparam ii3806.CONFIG_DATA = 16'h9A95;
      defparam ii3806.PLACE_LOCATION = "NONE";
      defparam ii3806.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3807 ( .DX(nn3807), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3763), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ) );
      defparam ii3807.CONFIG_DATA = 16'h9A95;
      defparam ii3807.PLACE_LOCATION = "NONE";
      defparam ii3807.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3808 ( .DX(nn3808), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3723), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ) );
      defparam ii3808.CONFIG_DATA = 16'h9A95;
      defparam ii3808.PLACE_LOCATION = "NONE";
      defparam ii3808.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3809 ( .DX(nn3809), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3725), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ) );
      defparam ii3809.CONFIG_DATA = 16'h9A95;
      defparam ii3809.PLACE_LOCATION = "NONE";
      defparam ii3809.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3810 ( .DX(nn3810), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3713), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_11|SUM_net ) );
      defparam ii3810.CONFIG_DATA = 16'h9A95;
      defparam ii3810.PLACE_LOCATION = "NONE";
      defparam ii3810.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3811 ( .DX(nn3811), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2694_), .F2(dummy_abc_2695_), .F3(dummy_abc_2696_) );
      defparam ii3811.CONFIG_DATA = 16'h5555;
      defparam ii3811.PLACE_LOCATION = "NONE";
      defparam ii3811.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3812 ( .DX(nn3812), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2697_), .F2(dummy_abc_2698_), .F3(dummy_abc_2699_) );
      defparam ii3812.CONFIG_DATA = 16'h5555;
      defparam ii3812.PLACE_LOCATION = "NONE";
      defparam ii3812.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3813 ( .DX(nn3813), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2700_), .F2(dummy_abc_2701_), .F3(dummy_abc_2702_) );
      defparam ii3813.CONFIG_DATA = 16'h5555;
      defparam ii3813.PLACE_LOCATION = "NONE";
      defparam ii3813.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3814 ( .DX(nn3814), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2703_), .F2(dummy_abc_2704_), .F3(dummy_abc_2705_) );
      defparam ii3814.CONFIG_DATA = 16'h5555;
      defparam ii3814.PLACE_LOCATION = "NONE";
      defparam ii3814.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3815 ( .DX(nn3815), .F0(dummy_abc_2706_), .F1(dummy_abc_2707_), .F2(dummy_abc_2708_), .F3(dummy_abc_2709_) );
      defparam ii3815.CONFIG_DATA = 16'hFFFF;
      defparam ii3815.PLACE_LOCATION = "NONE";
      defparam ii3815.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_240_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_432_ ), 
        .DX( {nn3815, nn3814, nn3813, nn3812, nn3811, nn3810, nn3809, nn3808, 
              nn3807, nn3806, nn3805, nn3804, nn3803, nn3802, nn3801, nn3800, 
              nn3755, nn3754} ), 
        .SUM( {\coefcal1_divide_inst1_u142_XORCI_17|SUM_net , dummy_433_, 
              dummy_434_, dummy_435_, dummy_436_, dummy_437_, dummy_438_, dummy_439_, 
              dummy_440_, dummy_441_, dummy_442_, dummy_443_, dummy_444_, dummy_445_, 
              dummy_446_, dummy_447_, dummy_448_, dummy_449_} )
      );
    CS_LUT4_PRIM ii3836 ( .DX(nn3836), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_413_), .F3(dummy_abc_2710_) );
      defparam ii3836.CONFIG_DATA = 16'hA6A6;
      defparam ii3836.PLACE_LOCATION = "NONE";
      defparam ii3836.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3837 ( .DX(nn3837), .F0(dummy_413_), .F1(nn3756), .F2(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ), .F3(dummy_abc_2711_) );
      defparam ii3837.CONFIG_DATA = 16'hD8D8;
      defparam ii3837.PLACE_LOCATION = "NONE";
      defparam ii3837.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3838 ( .DX(nn3838), .F0(nn3757), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ), .F3(dummy_abc_2712_) );
      defparam ii3838.CONFIG_DATA = 16'hB8B8;
      defparam ii3838.PLACE_LOCATION = "NONE";
      defparam ii3838.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3839 ( .DX(nn3839), .F0(nn3758), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ), .F3(dummy_abc_2713_) );
      defparam ii3839.CONFIG_DATA = 16'hB8B8;
      defparam ii3839.PLACE_LOCATION = "NONE";
      defparam ii3839.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3840 ( .DX(nn3840), .F0(nn3759), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ), .F3(dummy_abc_2714_) );
      defparam ii3840.CONFIG_DATA = 16'hB8B8;
      defparam ii3840.PLACE_LOCATION = "NONE";
      defparam ii3840.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3841 ( .DX(nn3841), .F0(nn3760), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ), .F3(dummy_abc_2715_) );
      defparam ii3841.CONFIG_DATA = 16'hB8B8;
      defparam ii3841.PLACE_LOCATION = "NONE";
      defparam ii3841.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3842 ( .DX(nn3842), .F0(nn3761), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ), .F3(dummy_abc_2716_) );
      defparam ii3842.CONFIG_DATA = 16'hB8B8;
      defparam ii3842.PLACE_LOCATION = "NONE";
      defparam ii3842.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3843 ( .DX(nn3843), .F0(nn3762), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ), .F3(dummy_abc_2717_) );
      defparam ii3843.CONFIG_DATA = 16'hB8B8;
      defparam ii3843.PLACE_LOCATION = "NONE";
      defparam ii3843.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3844 ( .DX(nn3844), .F0(nn3763), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ), .F3(dummy_abc_2718_) );
      defparam ii3844.CONFIG_DATA = 16'hB8B8;
      defparam ii3844.PLACE_LOCATION = "NONE";
      defparam ii3844.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3845 ( .DX(nn3845), .F0(nn3723), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ), .F3(dummy_abc_2719_) );
      defparam ii3845.CONFIG_DATA = 16'hB8B8;
      defparam ii3845.PLACE_LOCATION = "NONE";
      defparam ii3845.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3846 ( .DX(nn3846), .F0(nn3725), .F1(dummy_413_), .F2(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ), .F3(dummy_abc_2720_) );
      defparam ii3846.CONFIG_DATA = 16'hB8B8;
      defparam ii3846.PLACE_LOCATION = "NONE";
      defparam ii3846.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3847 ( .DX(nn3847), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2721_), .F3(dummy_abc_2722_) );
      defparam ii3847.CONFIG_DATA = 16'h9999;
      defparam ii3847.PLACE_LOCATION = "NONE";
      defparam ii3847.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3848 ( .DX(nn3848), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_413_) );
      defparam ii3848.CONFIG_DATA = 16'hA569;
      defparam ii3848.PLACE_LOCATION = "NONE";
      defparam ii3848.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3849 ( .DX(nn3849), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_413_), .F2(nn3756), .F3(\coefcal1_divide_inst1_u112_XORCI_1|SUM_net ) );
      defparam ii3849.CONFIG_DATA = 16'hA695;
      defparam ii3849.PLACE_LOCATION = "NONE";
      defparam ii3849.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3850 ( .DX(nn3850), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3757), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_2|SUM_net ) );
      defparam ii3850.CONFIG_DATA = 16'h9A95;
      defparam ii3850.PLACE_LOCATION = "NONE";
      defparam ii3850.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3851 ( .DX(nn3851), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3758), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_3|SUM_net ) );
      defparam ii3851.CONFIG_DATA = 16'h9A95;
      defparam ii3851.PLACE_LOCATION = "NONE";
      defparam ii3851.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3852 ( .DX(nn3852), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3759), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_4|SUM_net ) );
      defparam ii3852.CONFIG_DATA = 16'h9A95;
      defparam ii3852.PLACE_LOCATION = "NONE";
      defparam ii3852.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3853 ( .DX(nn3853), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3760), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_5|SUM_net ) );
      defparam ii3853.CONFIG_DATA = 16'h9A95;
      defparam ii3853.PLACE_LOCATION = "NONE";
      defparam ii3853.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3854 ( .DX(nn3854), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3761), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_6|SUM_net ) );
      defparam ii3854.CONFIG_DATA = 16'h9A95;
      defparam ii3854.PLACE_LOCATION = "NONE";
      defparam ii3854.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3855 ( .DX(nn3855), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3762), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_7|SUM_net ) );
      defparam ii3855.CONFIG_DATA = 16'h9A95;
      defparam ii3855.PLACE_LOCATION = "NONE";
      defparam ii3855.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3856 ( .DX(nn3856), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3763), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_8|SUM_net ) );
      defparam ii3856.CONFIG_DATA = 16'h9A95;
      defparam ii3856.PLACE_LOCATION = "NONE";
      defparam ii3856.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3857 ( .DX(nn3857), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3723), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_9|SUM_net ) );
      defparam ii3857.CONFIG_DATA = 16'h9A95;
      defparam ii3857.PLACE_LOCATION = "NONE";
      defparam ii3857.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3858 ( .DX(nn3858), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3725), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_10|SUM_net ) );
      defparam ii3858.CONFIG_DATA = 16'h9A95;
      defparam ii3858.PLACE_LOCATION = "NONE";
      defparam ii3858.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3859 ( .DX(nn3859), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3713), .F2(dummy_413_), .F3(\coefcal1_divide_inst1_u112_XORCI_11|SUM_net ) );
      defparam ii3859.CONFIG_DATA = 16'h9A95;
      defparam ii3859.PLACE_LOCATION = "NONE";
      defparam ii3859.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3860 ( .DX(nn3860), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(dummy_abc_2723_), .F2(dummy_abc_2724_), .F3(dummy_abc_2725_) );
      defparam ii3860.CONFIG_DATA = 16'h5555;
      defparam ii3860.PLACE_LOCATION = "NONE";
      defparam ii3860.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3861 ( .DX(nn3861), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2726_), .F2(dummy_abc_2727_), .F3(dummy_abc_2728_) );
      defparam ii3861.CONFIG_DATA = 16'h5555;
      defparam ii3861.PLACE_LOCATION = "NONE";
      defparam ii3861.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3862 ( .DX(nn3862), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2729_), .F2(dummy_abc_2730_), .F3(dummy_abc_2731_) );
      defparam ii3862.CONFIG_DATA = 16'h5555;
      defparam ii3862.PLACE_LOCATION = "NONE";
      defparam ii3862.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3863 ( .DX(nn3863), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2732_), .F2(dummy_abc_2733_), .F3(dummy_abc_2734_) );
      defparam ii3863.CONFIG_DATA = 16'h5555;
      defparam ii3863.PLACE_LOCATION = "NONE";
      defparam ii3863.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_225_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, nn3846, 
              nn3845, nn3844, nn3843, nn3842, nn3841, nn3840, nn3839, nn3838, 
              nn3837, nn3836, \coefcal1_xDividend__reg[4]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_163_ ), 
        .DX( {nn3863, nn3862, nn3861, nn3860, nn3859, nn3858, nn3857, nn3856, 
              nn3855, nn3854, nn3853, nn3852, nn3851, nn3850, nn3849, nn3848, 
              nn3847} ), 
        .SUM( {dummy_164_, \coefcal1_divide_inst1_u113_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_14|SUM_net , \coefcal1_divide_inst1_u113_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_12|SUM_net , \coefcal1_divide_inst1_u113_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_10|SUM_net , \coefcal1_divide_inst1_u113_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_8|SUM_net , \coefcal1_divide_inst1_u113_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_6|SUM_net , \coefcal1_divide_inst1_u113_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_4|SUM_net , \coefcal1_divide_inst1_u113_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_2|SUM_net , \coefcal1_divide_inst1_u113_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u113_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3883 ( .DX(nn3883), .F0(nn3713), .F1(dummy_413_), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3883.CONFIG_DATA = 16'h8F80;
      defparam ii3883.PLACE_LOCATION = "NONE";
      defparam ii3883.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3884 ( .DX(nn3884), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2735_), .F3(dummy_abc_2736_) );
      defparam ii3884.CONFIG_DATA = 16'h9999;
      defparam ii3884.PLACE_LOCATION = "NONE";
      defparam ii3884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3885 ( .DX(nn3885), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_432_) );
      defparam ii3885.CONFIG_DATA = 16'hA569;
      defparam ii3885.PLACE_LOCATION = "NONE";
      defparam ii3885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3886 ( .DX(nn3886), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_432_), .F2(nn3836), .F3(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ) );
      defparam ii3886.CONFIG_DATA = 16'hA695;
      defparam ii3886.PLACE_LOCATION = "NONE";
      defparam ii3886.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3887 ( .DX(nn3887), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3837), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ) );
      defparam ii3887.CONFIG_DATA = 16'h9A95;
      defparam ii3887.PLACE_LOCATION = "NONE";
      defparam ii3887.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3888 ( .DX(nn3888), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3838), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ) );
      defparam ii3888.CONFIG_DATA = 16'h9A95;
      defparam ii3888.PLACE_LOCATION = "NONE";
      defparam ii3888.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3889 ( .DX(nn3889), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3839), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ) );
      defparam ii3889.CONFIG_DATA = 16'h9A95;
      defparam ii3889.PLACE_LOCATION = "NONE";
      defparam ii3889.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3890 ( .DX(nn3890), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3840), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ) );
      defparam ii3890.CONFIG_DATA = 16'h9A95;
      defparam ii3890.PLACE_LOCATION = "NONE";
      defparam ii3890.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3891 ( .DX(nn3891), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3841), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ) );
      defparam ii3891.CONFIG_DATA = 16'h9A95;
      defparam ii3891.PLACE_LOCATION = "NONE";
      defparam ii3891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3892 ( .DX(nn3892), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3842), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ) );
      defparam ii3892.CONFIG_DATA = 16'h9A95;
      defparam ii3892.PLACE_LOCATION = "NONE";
      defparam ii3892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3893 ( .DX(nn3893), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3843), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ) );
      defparam ii3893.CONFIG_DATA = 16'h9A95;
      defparam ii3893.PLACE_LOCATION = "NONE";
      defparam ii3893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3894 ( .DX(nn3894), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3844), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ) );
      defparam ii3894.CONFIG_DATA = 16'h9A95;
      defparam ii3894.PLACE_LOCATION = "NONE";
      defparam ii3894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3895 ( .DX(nn3895), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3845), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ) );
      defparam ii3895.CONFIG_DATA = 16'h9A95;
      defparam ii3895.PLACE_LOCATION = "NONE";
      defparam ii3895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3896 ( .DX(nn3896), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3846), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ) );
      defparam ii3896.CONFIG_DATA = 16'h9A95;
      defparam ii3896.PLACE_LOCATION = "NONE";
      defparam ii3896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3897 ( .DX(nn3897), .F0(nn3713), .F1(dummy_413_), .F2(dummy_abc_2737_), .F3(dummy_abc_2738_) );
      defparam ii3897.CONFIG_DATA = 16'h8888;
      defparam ii3897.PLACE_LOCATION = "NONE";
      defparam ii3897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3898 ( .DX(nn3898), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3897), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3898.CONFIG_DATA = 16'h9095;
      defparam ii3898.PLACE_LOCATION = "NONE";
      defparam ii3898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3899 ( .DX(nn3899), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2739_), .F2(dummy_abc_2740_), .F3(dummy_abc_2741_) );
      defparam ii3899.CONFIG_DATA = 16'h5555;
      defparam ii3899.PLACE_LOCATION = "NONE";
      defparam ii3899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3900 ( .DX(nn3900), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2742_), .F2(dummy_abc_2743_), .F3(dummy_abc_2744_) );
      defparam ii3900.CONFIG_DATA = 16'h5555;
      defparam ii3900.PLACE_LOCATION = "NONE";
      defparam ii3900.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3901 ( .DX(nn3901), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2745_), .F2(dummy_abc_2746_), .F3(dummy_abc_2747_) );
      defparam ii3901.CONFIG_DATA = 16'h5555;
      defparam ii3901.PLACE_LOCATION = "NONE";
      defparam ii3901.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3902 ( .DX(nn3902), .F0(dummy_abc_2748_), .F1(dummy_abc_2749_), .F2(dummy_abc_2750_), .F3(dummy_abc_2751_) );
      defparam ii3902.CONFIG_DATA = 16'hFFFF;
      defparam ii3902.PLACE_LOCATION = "NONE";
      defparam ii3902.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_241_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_451_ ), 
        .DX( {nn3902, nn3901, nn3900, nn3899, nn3898, nn3896, nn3895, nn3894, 
              nn3893, nn3892, nn3891, nn3890, nn3889, nn3888, nn3887, nn3886, 
              nn3885, nn3884} ), 
        .SUM( {\coefcal1_divide_inst1_u144_XORCI_17|SUM_net , dummy_452_, 
              dummy_453_, dummy_454_, dummy_455_, dummy_456_, dummy_457_, dummy_458_, 
              dummy_459_, dummy_460_, dummy_461_, dummy_462_, dummy_463_, dummy_464_, 
              dummy_465_, dummy_466_, dummy_467_, dummy_468_} )
      );
    CS_LUT4_PRIM ii3923 ( .DX(nn3923), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_432_), .F3(dummy_abc_2752_) );
      defparam ii3923.CONFIG_DATA = 16'hA6A6;
      defparam ii3923.PLACE_LOCATION = "NONE";
      defparam ii3923.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3924 ( .DX(nn3924), .F0(dummy_432_), .F1(nn3836), .F2(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ), .F3(dummy_abc_2753_) );
      defparam ii3924.CONFIG_DATA = 16'hD8D8;
      defparam ii3924.PLACE_LOCATION = "NONE";
      defparam ii3924.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3925 ( .DX(nn3925), .F0(nn3837), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ), .F3(dummy_abc_2754_) );
      defparam ii3925.CONFIG_DATA = 16'hB8B8;
      defparam ii3925.PLACE_LOCATION = "NONE";
      defparam ii3925.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3926 ( .DX(nn3926), .F0(nn3838), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ), .F3(dummy_abc_2755_) );
      defparam ii3926.CONFIG_DATA = 16'hB8B8;
      defparam ii3926.PLACE_LOCATION = "NONE";
      defparam ii3926.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3927 ( .DX(nn3927), .F0(nn3839), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ), .F3(dummy_abc_2756_) );
      defparam ii3927.CONFIG_DATA = 16'hB8B8;
      defparam ii3927.PLACE_LOCATION = "NONE";
      defparam ii3927.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3928 ( .DX(nn3928), .F0(nn3840), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ), .F3(dummy_abc_2757_) );
      defparam ii3928.CONFIG_DATA = 16'hB8B8;
      defparam ii3928.PLACE_LOCATION = "NONE";
      defparam ii3928.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3929 ( .DX(nn3929), .F0(nn3841), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ), .F3(dummy_abc_2758_) );
      defparam ii3929.CONFIG_DATA = 16'hB8B8;
      defparam ii3929.PLACE_LOCATION = "NONE";
      defparam ii3929.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3930 ( .DX(nn3930), .F0(nn3842), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ), .F3(dummy_abc_2759_) );
      defparam ii3930.CONFIG_DATA = 16'hB8B8;
      defparam ii3930.PLACE_LOCATION = "NONE";
      defparam ii3930.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3931 ( .DX(nn3931), .F0(nn3843), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ), .F3(dummy_abc_2760_) );
      defparam ii3931.CONFIG_DATA = 16'hB8B8;
      defparam ii3931.PLACE_LOCATION = "NONE";
      defparam ii3931.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3932 ( .DX(nn3932), .F0(nn3844), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ), .F3(dummy_abc_2761_) );
      defparam ii3932.CONFIG_DATA = 16'hB8B8;
      defparam ii3932.PLACE_LOCATION = "NONE";
      defparam ii3932.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3933 ( .DX(nn3933), .F0(nn3845), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ), .F3(dummy_abc_2762_) );
      defparam ii3933.CONFIG_DATA = 16'hB8B8;
      defparam ii3933.PLACE_LOCATION = "NONE";
      defparam ii3933.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3934 ( .DX(nn3934), .F0(nn3846), .F1(dummy_432_), .F2(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ), .F3(dummy_abc_2763_) );
      defparam ii3934.CONFIG_DATA = 16'hB8B8;
      defparam ii3934.PLACE_LOCATION = "NONE";
      defparam ii3934.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3935 ( .DX(nn3935), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2764_), .F3(dummy_abc_2765_) );
      defparam ii3935.CONFIG_DATA = 16'h9999;
      defparam ii3935.PLACE_LOCATION = "NONE";
      defparam ii3935.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3936 ( .DX(nn3936), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_432_) );
      defparam ii3936.CONFIG_DATA = 16'hA569;
      defparam ii3936.PLACE_LOCATION = "NONE";
      defparam ii3936.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3937 ( .DX(nn3937), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_432_), .F2(nn3836), .F3(\coefcal1_divide_inst1_u113_XORCI_1|SUM_net ) );
      defparam ii3937.CONFIG_DATA = 16'hA695;
      defparam ii3937.PLACE_LOCATION = "NONE";
      defparam ii3937.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3938 ( .DX(nn3938), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3837), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_2|SUM_net ) );
      defparam ii3938.CONFIG_DATA = 16'h9A95;
      defparam ii3938.PLACE_LOCATION = "NONE";
      defparam ii3938.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3939 ( .DX(nn3939), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3838), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_3|SUM_net ) );
      defparam ii3939.CONFIG_DATA = 16'h9A95;
      defparam ii3939.PLACE_LOCATION = "NONE";
      defparam ii3939.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3940 ( .DX(nn3940), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3839), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_4|SUM_net ) );
      defparam ii3940.CONFIG_DATA = 16'h9A95;
      defparam ii3940.PLACE_LOCATION = "NONE";
      defparam ii3940.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3941 ( .DX(nn3941), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3840), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_5|SUM_net ) );
      defparam ii3941.CONFIG_DATA = 16'h9A95;
      defparam ii3941.PLACE_LOCATION = "NONE";
      defparam ii3941.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3942 ( .DX(nn3942), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3841), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_6|SUM_net ) );
      defparam ii3942.CONFIG_DATA = 16'h9A95;
      defparam ii3942.PLACE_LOCATION = "NONE";
      defparam ii3942.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3943 ( .DX(nn3943), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3842), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_7|SUM_net ) );
      defparam ii3943.CONFIG_DATA = 16'h9A95;
      defparam ii3943.PLACE_LOCATION = "NONE";
      defparam ii3943.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3944 ( .DX(nn3944), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3843), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_8|SUM_net ) );
      defparam ii3944.CONFIG_DATA = 16'h9A95;
      defparam ii3944.PLACE_LOCATION = "NONE";
      defparam ii3944.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3945 ( .DX(nn3945), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3844), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_9|SUM_net ) );
      defparam ii3945.CONFIG_DATA = 16'h9A95;
      defparam ii3945.PLACE_LOCATION = "NONE";
      defparam ii3945.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3946 ( .DX(nn3946), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3845), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_10|SUM_net ) );
      defparam ii3946.CONFIG_DATA = 16'h9A95;
      defparam ii3946.PLACE_LOCATION = "NONE";
      defparam ii3946.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3947 ( .DX(nn3947), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3846), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_11|SUM_net ) );
      defparam ii3947.CONFIG_DATA = 16'h9A95;
      defparam ii3947.PLACE_LOCATION = "NONE";
      defparam ii3947.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3948 ( .DX(nn3948), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3897), .F2(dummy_432_), .F3(\coefcal1_divide_inst1_u113_XORCI_12|SUM_net ) );
      defparam ii3948.CONFIG_DATA = 16'h9095;
      defparam ii3948.PLACE_LOCATION = "NONE";
      defparam ii3948.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3949 ( .DX(nn3949), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(dummy_abc_2766_), .F2(dummy_abc_2767_), .F3(dummy_abc_2768_) );
      defparam ii3949.CONFIG_DATA = 16'h5555;
      defparam ii3949.PLACE_LOCATION = "NONE";
      defparam ii3949.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3950 ( .DX(nn3950), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2769_), .F2(dummy_abc_2770_), .F3(dummy_abc_2771_) );
      defparam ii3950.CONFIG_DATA = 16'h5555;
      defparam ii3950.PLACE_LOCATION = "NONE";
      defparam ii3950.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3951 ( .DX(nn3951), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2772_), .F2(dummy_abc_2773_), .F3(dummy_abc_2774_) );
      defparam ii3951.CONFIG_DATA = 16'h5555;
      defparam ii3951.PLACE_LOCATION = "NONE";
      defparam ii3951.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_226_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn3883, nn3934, nn3933, nn3932, nn3931, nn3930, nn3929, 
              nn3928, nn3927, nn3926, nn3925, nn3924, nn3923, 
              \coefcal1_xDividend__reg[3]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_165_ ), 
        .DX( {nn3951, nn3950, nn3949, nn3948, nn3947, nn3946, nn3945, nn3944, 
              nn3943, nn3942, nn3941, nn3940, nn3939, nn3938, nn3937, nn3936, 
              nn3935} ), 
        .SUM( {dummy_166_, \coefcal1_divide_inst1_u114_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_14|SUM_net , \coefcal1_divide_inst1_u114_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_12|SUM_net , \coefcal1_divide_inst1_u114_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_10|SUM_net , \coefcal1_divide_inst1_u114_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_8|SUM_net , \coefcal1_divide_inst1_u114_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_6|SUM_net , \coefcal1_divide_inst1_u114_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_4|SUM_net , \coefcal1_divide_inst1_u114_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_2|SUM_net , \coefcal1_divide_inst1_u114_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u114_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii3971 ( .DX(nn3971), .F0(dummy_451_), .F1(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ), .F2(dummy_abc_2775_), .F3(dummy_abc_2776_) );
      defparam ii3971.CONFIG_DATA = 16'h1111;
      defparam ii3971.PLACE_LOCATION = "NONE";
      defparam ii3971.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3972 ( .DX(nn3972), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2777_), .F3(dummy_abc_2778_) );
      defparam ii3972.CONFIG_DATA = 16'h9999;
      defparam ii3972.PLACE_LOCATION = "NONE";
      defparam ii3972.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3973 ( .DX(nn3973), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_451_) );
      defparam ii3973.CONFIG_DATA = 16'hA569;
      defparam ii3973.PLACE_LOCATION = "NONE";
      defparam ii3973.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3974 ( .DX(nn3974), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_451_), .F2(nn3923), .F3(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ) );
      defparam ii3974.CONFIG_DATA = 16'hA695;
      defparam ii3974.PLACE_LOCATION = "NONE";
      defparam ii3974.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3975 ( .DX(nn3975), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3924), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ) );
      defparam ii3975.CONFIG_DATA = 16'h9A95;
      defparam ii3975.PLACE_LOCATION = "NONE";
      defparam ii3975.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3976 ( .DX(nn3976), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3925), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ) );
      defparam ii3976.CONFIG_DATA = 16'h9A95;
      defparam ii3976.PLACE_LOCATION = "NONE";
      defparam ii3976.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3977 ( .DX(nn3977), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3926), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ) );
      defparam ii3977.CONFIG_DATA = 16'h9A95;
      defparam ii3977.PLACE_LOCATION = "NONE";
      defparam ii3977.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3978 ( .DX(nn3978), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3927), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ) );
      defparam ii3978.CONFIG_DATA = 16'h9A95;
      defparam ii3978.PLACE_LOCATION = "NONE";
      defparam ii3978.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3979 ( .DX(nn3979), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3928), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ) );
      defparam ii3979.CONFIG_DATA = 16'h9A95;
      defparam ii3979.PLACE_LOCATION = "NONE";
      defparam ii3979.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3980 ( .DX(nn3980), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3929), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ) );
      defparam ii3980.CONFIG_DATA = 16'h9A95;
      defparam ii3980.PLACE_LOCATION = "NONE";
      defparam ii3980.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3981 ( .DX(nn3981), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3930), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ) );
      defparam ii3981.CONFIG_DATA = 16'h9A95;
      defparam ii3981.PLACE_LOCATION = "NONE";
      defparam ii3981.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3982 ( .DX(nn3982), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3931), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ) );
      defparam ii3982.CONFIG_DATA = 16'h9A95;
      defparam ii3982.PLACE_LOCATION = "NONE";
      defparam ii3982.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3983 ( .DX(nn3983), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3932), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ) );
      defparam ii3983.CONFIG_DATA = 16'h9A95;
      defparam ii3983.PLACE_LOCATION = "NONE";
      defparam ii3983.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3984 ( .DX(nn3984), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3933), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ) );
      defparam ii3984.CONFIG_DATA = 16'h9A95;
      defparam ii3984.PLACE_LOCATION = "NONE";
      defparam ii3984.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3985 ( .DX(nn3985), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3934), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ) );
      defparam ii3985.CONFIG_DATA = 16'h9A95;
      defparam ii3985.PLACE_LOCATION = "NONE";
      defparam ii3985.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3986 ( .DX(nn3986), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3883), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ) );
      defparam ii3986.CONFIG_DATA = 16'h9995;
      defparam ii3986.PLACE_LOCATION = "NONE";
      defparam ii3986.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3987 ( .DX(nn3987), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2779_), .F2(dummy_abc_2780_), .F3(dummy_abc_2781_) );
      defparam ii3987.CONFIG_DATA = 16'h5555;
      defparam ii3987.PLACE_LOCATION = "NONE";
      defparam ii3987.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3988 ( .DX(nn3988), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2782_), .F2(dummy_abc_2783_), .F3(dummy_abc_2784_) );
      defparam ii3988.CONFIG_DATA = 16'h5555;
      defparam ii3988.PLACE_LOCATION = "NONE";
      defparam ii3988.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii3989 ( .DX(nn3989), .F0(dummy_abc_2785_), .F1(dummy_abc_2786_), .F2(dummy_abc_2787_), .F3(dummy_abc_2788_) );
      defparam ii3989.CONFIG_DATA = 16'hFFFF;
      defparam ii3989.PLACE_LOCATION = "NONE";
      defparam ii3989.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_242_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_470_ ), 
        .DX( {nn3989, nn3988, nn3987, nn3986, nn3985, nn3984, nn3983, nn3982, 
              nn3981, nn3980, nn3979, nn3978, nn3977, nn3976, nn3975, nn3974, 
              nn3973, nn3972} ), 
        .SUM( {\coefcal1_divide_inst1_u146_XORCI_17|SUM_net , dummy_471_, 
              dummy_472_, dummy_473_, dummy_474_, dummy_475_, dummy_476_, dummy_477_, 
              dummy_478_, dummy_479_, dummy_480_, dummy_481_, dummy_482_, dummy_483_, 
              dummy_484_, dummy_485_, dummy_486_, dummy_487_} )
      );
    CS_LUT4_PRIM ii4010 ( .DX(nn4010), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_451_), .F3(dummy_abc_2789_) );
      defparam ii4010.CONFIG_DATA = 16'hA6A6;
      defparam ii4010.PLACE_LOCATION = "NONE";
      defparam ii4010.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4011 ( .DX(nn4011), .F0(dummy_451_), .F1(nn3923), .F2(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ), .F3(dummy_abc_2790_) );
      defparam ii4011.CONFIG_DATA = 16'hD8D8;
      defparam ii4011.PLACE_LOCATION = "NONE";
      defparam ii4011.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4012 ( .DX(nn4012), .F0(nn3924), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ), .F3(dummy_abc_2791_) );
      defparam ii4012.CONFIG_DATA = 16'hB8B8;
      defparam ii4012.PLACE_LOCATION = "NONE";
      defparam ii4012.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4013 ( .DX(nn4013), .F0(nn3925), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ), .F3(dummy_abc_2792_) );
      defparam ii4013.CONFIG_DATA = 16'hB8B8;
      defparam ii4013.PLACE_LOCATION = "NONE";
      defparam ii4013.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4014 ( .DX(nn4014), .F0(nn3926), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ), .F3(dummy_abc_2793_) );
      defparam ii4014.CONFIG_DATA = 16'hB8B8;
      defparam ii4014.PLACE_LOCATION = "NONE";
      defparam ii4014.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4015 ( .DX(nn4015), .F0(nn3927), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ), .F3(dummy_abc_2794_) );
      defparam ii4015.CONFIG_DATA = 16'hB8B8;
      defparam ii4015.PLACE_LOCATION = "NONE";
      defparam ii4015.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4016 ( .DX(nn4016), .F0(nn3928), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ), .F3(dummy_abc_2795_) );
      defparam ii4016.CONFIG_DATA = 16'hB8B8;
      defparam ii4016.PLACE_LOCATION = "NONE";
      defparam ii4016.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4017 ( .DX(nn4017), .F0(nn3929), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ), .F3(dummy_abc_2796_) );
      defparam ii4017.CONFIG_DATA = 16'hB8B8;
      defparam ii4017.PLACE_LOCATION = "NONE";
      defparam ii4017.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4018 ( .DX(nn4018), .F0(nn3930), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ), .F3(dummy_abc_2797_) );
      defparam ii4018.CONFIG_DATA = 16'hB8B8;
      defparam ii4018.PLACE_LOCATION = "NONE";
      defparam ii4018.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4019 ( .DX(nn4019), .F0(nn3931), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ), .F3(dummy_abc_2798_) );
      defparam ii4019.CONFIG_DATA = 16'hB8B8;
      defparam ii4019.PLACE_LOCATION = "NONE";
      defparam ii4019.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4020 ( .DX(nn4020), .F0(nn3932), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ), .F3(dummy_abc_2799_) );
      defparam ii4020.CONFIG_DATA = 16'hB8B8;
      defparam ii4020.PLACE_LOCATION = "NONE";
      defparam ii4020.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4021 ( .DX(nn4021), .F0(nn3933), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ), .F3(dummy_abc_2800_) );
      defparam ii4021.CONFIG_DATA = 16'hB8B8;
      defparam ii4021.PLACE_LOCATION = "NONE";
      defparam ii4021.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4022 ( .DX(nn4022), .F0(nn3934), .F1(dummy_451_), .F2(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ), .F3(dummy_abc_2801_) );
      defparam ii4022.CONFIG_DATA = 16'hB8B8;
      defparam ii4022.PLACE_LOCATION = "NONE";
      defparam ii4022.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4023 ( .DX(nn4023), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2802_), .F3(dummy_abc_2803_) );
      defparam ii4023.CONFIG_DATA = 16'h9999;
      defparam ii4023.PLACE_LOCATION = "NONE";
      defparam ii4023.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4024 ( .DX(nn4024), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_451_) );
      defparam ii4024.CONFIG_DATA = 16'hA569;
      defparam ii4024.PLACE_LOCATION = "NONE";
      defparam ii4024.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4025 ( .DX(nn4025), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_451_), .F2(nn3923), .F3(\coefcal1_divide_inst1_u114_XORCI_1|SUM_net ) );
      defparam ii4025.CONFIG_DATA = 16'hA695;
      defparam ii4025.PLACE_LOCATION = "NONE";
      defparam ii4025.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4026 ( .DX(nn4026), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn3924), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_2|SUM_net ) );
      defparam ii4026.CONFIG_DATA = 16'h9A95;
      defparam ii4026.PLACE_LOCATION = "NONE";
      defparam ii4026.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4027 ( .DX(nn4027), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn3925), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_3|SUM_net ) );
      defparam ii4027.CONFIG_DATA = 16'h9A95;
      defparam ii4027.PLACE_LOCATION = "NONE";
      defparam ii4027.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4028 ( .DX(nn4028), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn3926), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_4|SUM_net ) );
      defparam ii4028.CONFIG_DATA = 16'h9A95;
      defparam ii4028.PLACE_LOCATION = "NONE";
      defparam ii4028.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4029 ( .DX(nn4029), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn3927), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_5|SUM_net ) );
      defparam ii4029.CONFIG_DATA = 16'h9A95;
      defparam ii4029.PLACE_LOCATION = "NONE";
      defparam ii4029.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4030 ( .DX(nn4030), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn3928), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_6|SUM_net ) );
      defparam ii4030.CONFIG_DATA = 16'h9A95;
      defparam ii4030.PLACE_LOCATION = "NONE";
      defparam ii4030.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4031 ( .DX(nn4031), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn3929), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_7|SUM_net ) );
      defparam ii4031.CONFIG_DATA = 16'h9A95;
      defparam ii4031.PLACE_LOCATION = "NONE";
      defparam ii4031.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4032 ( .DX(nn4032), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn3930), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_8|SUM_net ) );
      defparam ii4032.CONFIG_DATA = 16'h9A95;
      defparam ii4032.PLACE_LOCATION = "NONE";
      defparam ii4032.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4033 ( .DX(nn4033), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn3931), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_9|SUM_net ) );
      defparam ii4033.CONFIG_DATA = 16'h9A95;
      defparam ii4033.PLACE_LOCATION = "NONE";
      defparam ii4033.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4034 ( .DX(nn4034), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn3932), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_10|SUM_net ) );
      defparam ii4034.CONFIG_DATA = 16'h9A95;
      defparam ii4034.PLACE_LOCATION = "NONE";
      defparam ii4034.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4035 ( .DX(nn4035), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn3933), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_11|SUM_net ) );
      defparam ii4035.CONFIG_DATA = 16'h9A95;
      defparam ii4035.PLACE_LOCATION = "NONE";
      defparam ii4035.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4036 ( .DX(nn4036), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn3934), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_12|SUM_net ) );
      defparam ii4036.CONFIG_DATA = 16'h9A95;
      defparam ii4036.PLACE_LOCATION = "NONE";
      defparam ii4036.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4037 ( .DX(nn4037), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn3883), .F2(dummy_451_), .F3(\coefcal1_divide_inst1_u114_XORCI_13|SUM_net ) );
      defparam ii4037.CONFIG_DATA = 16'h9995;
      defparam ii4037.PLACE_LOCATION = "NONE";
      defparam ii4037.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4038 ( .DX(nn4038), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(dummy_abc_2804_), .F2(dummy_abc_2805_), .F3(dummy_abc_2806_) );
      defparam ii4038.CONFIG_DATA = 16'h5555;
      defparam ii4038.PLACE_LOCATION = "NONE";
      defparam ii4038.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4039 ( .DX(nn4039), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2807_), .F2(dummy_abc_2808_), .F3(dummy_abc_2809_) );
      defparam ii4039.CONFIG_DATA = 16'h5555;
      defparam ii4039.PLACE_LOCATION = "NONE";
      defparam ii4039.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_227_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, nn4022, nn4021, nn4020, nn4019, nn4018, nn4017, nn4016, 
              nn4015, nn4014, nn4013, nn4012, nn4011, nn4010, 
              \coefcal1_xDividend__reg[2]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_167_ ), 
        .DX( {nn4039, nn4038, nn4037, nn4036, nn4035, nn4034, nn4033, nn4032, 
              nn4031, nn4030, nn4029, nn4028, nn4027, nn4026, nn4025, nn4024, 
              nn4023} ), 
        .SUM( {dummy_168_, \coefcal1_divide_inst1_u115_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_14|SUM_net , \coefcal1_divide_inst1_u115_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_12|SUM_net , \coefcal1_divide_inst1_u115_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_10|SUM_net , \coefcal1_divide_inst1_u115_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_8|SUM_net , \coefcal1_divide_inst1_u115_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_6|SUM_net , \coefcal1_divide_inst1_u115_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_4|SUM_net , \coefcal1_divide_inst1_u115_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_2|SUM_net , \coefcal1_divide_inst1_u115_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u115_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4059 ( .DX(nn4059), .F0(nn3883), .F1(nn3971), .F2(dummy_470_), .F3(\coefcal1_divide_inst1_u115_XORCI_14|SUM_net ) );
      defparam ii4059.CONFIG_DATA = 16'h2A20;
      defparam ii4059.PLACE_LOCATION = "NONE";
      defparam ii4059.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4060 ( .DX(nn4060), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2810_), .F3(dummy_abc_2811_) );
      defparam ii4060.CONFIG_DATA = 16'h9999;
      defparam ii4060.PLACE_LOCATION = "NONE";
      defparam ii4060.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4061 ( .DX(nn4061), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_470_) );
      defparam ii4061.CONFIG_DATA = 16'hA569;
      defparam ii4061.PLACE_LOCATION = "NONE";
      defparam ii4061.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4062 ( .DX(nn4062), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_470_), .F2(nn4010), .F3(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ) );
      defparam ii4062.CONFIG_DATA = 16'hA695;
      defparam ii4062.PLACE_LOCATION = "NONE";
      defparam ii4062.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4063 ( .DX(nn4063), .F0(nn4011), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_2|SUM_net ), .F3(dummy_abc_2812_) );
      defparam ii4063.CONFIG_DATA = 16'hB8B8;
      defparam ii4063.PLACE_LOCATION = "NONE";
      defparam ii4063.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4064 ( .DX(nn4064), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn4063), .F2(dummy_abc_2813_), .F3(dummy_abc_2814_) );
      defparam ii4064.CONFIG_DATA = 16'h9999;
      defparam ii4064.PLACE_LOCATION = "NONE";
      defparam ii4064.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4065 ( .DX(nn4065), .F0(nn4012), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_3|SUM_net ), .F3(dummy_abc_2815_) );
      defparam ii4065.CONFIG_DATA = 16'hB8B8;
      defparam ii4065.PLACE_LOCATION = "NONE";
      defparam ii4065.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4066 ( .DX(nn4066), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn4065), .F2(dummy_abc_2816_), .F3(dummy_abc_2817_) );
      defparam ii4066.CONFIG_DATA = 16'h9999;
      defparam ii4066.PLACE_LOCATION = "NONE";
      defparam ii4066.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4067 ( .DX(nn4067), .F0(nn4013), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_4|SUM_net ), .F3(dummy_abc_2818_) );
      defparam ii4067.CONFIG_DATA = 16'hB8B8;
      defparam ii4067.PLACE_LOCATION = "NONE";
      defparam ii4067.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4068 ( .DX(nn4068), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn4067), .F2(dummy_abc_2819_), .F3(dummy_abc_2820_) );
      defparam ii4068.CONFIG_DATA = 16'h9999;
      defparam ii4068.PLACE_LOCATION = "NONE";
      defparam ii4068.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4069 ( .DX(nn4069), .F0(nn4014), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_5|SUM_net ), .F3(dummy_abc_2821_) );
      defparam ii4069.CONFIG_DATA = 16'hB8B8;
      defparam ii4069.PLACE_LOCATION = "NONE";
      defparam ii4069.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4070 ( .DX(nn4070), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn4069), .F2(dummy_abc_2822_), .F3(dummy_abc_2823_) );
      defparam ii4070.CONFIG_DATA = 16'h9999;
      defparam ii4070.PLACE_LOCATION = "NONE";
      defparam ii4070.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4071 ( .DX(nn4071), .F0(nn4015), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_6|SUM_net ), .F3(dummy_abc_2824_) );
      defparam ii4071.CONFIG_DATA = 16'hB8B8;
      defparam ii4071.PLACE_LOCATION = "NONE";
      defparam ii4071.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4072 ( .DX(nn4072), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn4071), .F2(dummy_abc_2825_), .F3(dummy_abc_2826_) );
      defparam ii4072.CONFIG_DATA = 16'h9999;
      defparam ii4072.PLACE_LOCATION = "NONE";
      defparam ii4072.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4073 ( .DX(nn4073), .F0(nn4016), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_7|SUM_net ), .F3(dummy_abc_2827_) );
      defparam ii4073.CONFIG_DATA = 16'hB8B8;
      defparam ii4073.PLACE_LOCATION = "NONE";
      defparam ii4073.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4074 ( .DX(nn4074), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn4073), .F2(dummy_abc_2828_), .F3(dummy_abc_2829_) );
      defparam ii4074.CONFIG_DATA = 16'h9999;
      defparam ii4074.PLACE_LOCATION = "NONE";
      defparam ii4074.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4075 ( .DX(nn4075), .F0(nn4017), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_8|SUM_net ), .F3(dummy_abc_2830_) );
      defparam ii4075.CONFIG_DATA = 16'hB8B8;
      defparam ii4075.PLACE_LOCATION = "NONE";
      defparam ii4075.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4076 ( .DX(nn4076), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn4075), .F2(dummy_abc_2831_), .F3(dummy_abc_2832_) );
      defparam ii4076.CONFIG_DATA = 16'h9999;
      defparam ii4076.PLACE_LOCATION = "NONE";
      defparam ii4076.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4077 ( .DX(nn4077), .F0(nn4018), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_9|SUM_net ), .F3(dummy_abc_2833_) );
      defparam ii4077.CONFIG_DATA = 16'hB8B8;
      defparam ii4077.PLACE_LOCATION = "NONE";
      defparam ii4077.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4078 ( .DX(nn4078), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn4077), .F2(dummy_abc_2834_), .F3(dummy_abc_2835_) );
      defparam ii4078.CONFIG_DATA = 16'h9999;
      defparam ii4078.PLACE_LOCATION = "NONE";
      defparam ii4078.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4079 ( .DX(nn4079), .F0(nn4019), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_10|SUM_net ), .F3(dummy_abc_2836_) );
      defparam ii4079.CONFIG_DATA = 16'hB8B8;
      defparam ii4079.PLACE_LOCATION = "NONE";
      defparam ii4079.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4080 ( .DX(nn4080), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn4079), .F2(dummy_abc_2837_), .F3(dummy_abc_2838_) );
      defparam ii4080.CONFIG_DATA = 16'h9999;
      defparam ii4080.PLACE_LOCATION = "NONE";
      defparam ii4080.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4081 ( .DX(nn4081), .F0(nn4020), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_11|SUM_net ), .F3(dummy_abc_2839_) );
      defparam ii4081.CONFIG_DATA = 16'hB8B8;
      defparam ii4081.PLACE_LOCATION = "NONE";
      defparam ii4081.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4082 ( .DX(nn4082), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn4081), .F2(dummy_abc_2840_), .F3(dummy_abc_2841_) );
      defparam ii4082.CONFIG_DATA = 16'h9999;
      defparam ii4082.PLACE_LOCATION = "NONE";
      defparam ii4082.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4083 ( .DX(nn4083), .F0(nn4021), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_12|SUM_net ), .F3(dummy_abc_2842_) );
      defparam ii4083.CONFIG_DATA = 16'hB8B8;
      defparam ii4083.PLACE_LOCATION = "NONE";
      defparam ii4083.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4084 ( .DX(nn4084), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn4083), .F2(dummy_abc_2843_), .F3(dummy_abc_2844_) );
      defparam ii4084.CONFIG_DATA = 16'h9999;
      defparam ii4084.PLACE_LOCATION = "NONE";
      defparam ii4084.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4085 ( .DX(nn4085), .F0(nn4022), .F1(dummy_470_), .F2(\coefcal1_divide_inst1_u115_XORCI_13|SUM_net ), .F3(dummy_abc_2845_) );
      defparam ii4085.CONFIG_DATA = 16'hB8B8;
      defparam ii4085.PLACE_LOCATION = "NONE";
      defparam ii4085.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4086 ( .DX(nn4086), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn4085), .F2(dummy_abc_2846_), .F3(dummy_abc_2847_) );
      defparam ii4086.CONFIG_DATA = 16'h9999;
      defparam ii4086.PLACE_LOCATION = "NONE";
      defparam ii4086.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4087 ( .DX(nn4087), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn4059), .F2(dummy_abc_2848_), .F3(dummy_abc_2849_) );
      defparam ii4087.CONFIG_DATA = 16'h9999;
      defparam ii4087.PLACE_LOCATION = "NONE";
      defparam ii4087.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4088 ( .DX(nn4088), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2850_), .F2(dummy_abc_2851_), .F3(dummy_abc_2852_) );
      defparam ii4088.CONFIG_DATA = 16'h5555;
      defparam ii4088.PLACE_LOCATION = "NONE";
      defparam ii4088.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4089 ( .DX(nn4089), .F0(dummy_abc_2853_), .F1(dummy_abc_2854_), .F2(dummy_abc_2855_), .F3(dummy_abc_2856_) );
      defparam ii4089.CONFIG_DATA = 16'hFFFF;
      defparam ii4089.PLACE_LOCATION = "NONE";
      defparam ii4089.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_243_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_489_ ), 
        .DX( {nn4089, nn4088, nn4087, nn4086, nn4084, nn4082, nn4080, nn4078, 
              nn4076, nn4074, nn4072, nn4070, nn4068, nn4066, nn4064, nn4062, 
              nn4061, nn4060} ), 
        .SUM( {\coefcal1_divide_inst1_u148_XORCI_17|SUM_net , dummy_490_, 
              dummy_491_, dummy_492_, dummy_493_, dummy_494_, dummy_495_, dummy_496_, 
              dummy_497_, dummy_498_, dummy_499_, dummy_500_, dummy_501_, dummy_502_, 
              dummy_503_, dummy_504_, dummy_505_, dummy_506_} )
      );
    CS_LUT4_PRIM ii4110 ( .DX(nn4110), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_470_), .F3(dummy_abc_2857_) );
      defparam ii4110.CONFIG_DATA = 16'hA6A6;
      defparam ii4110.PLACE_LOCATION = "NONE";
      defparam ii4110.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4111 ( .DX(nn4111), .F0(dummy_470_), .F1(nn4010), .F2(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ), .F3(dummy_abc_2858_) );
      defparam ii4111.CONFIG_DATA = 16'hD8D8;
      defparam ii4111.PLACE_LOCATION = "NONE";
      defparam ii4111.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4112 ( .DX(nn4112), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2859_), .F3(dummy_abc_2860_) );
      defparam ii4112.CONFIG_DATA = 16'h9999;
      defparam ii4112.PLACE_LOCATION = "NONE";
      defparam ii4112.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4113 ( .DX(nn4113), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_470_) );
      defparam ii4113.CONFIG_DATA = 16'hA569;
      defparam ii4113.PLACE_LOCATION = "NONE";
      defparam ii4113.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4114 ( .DX(nn4114), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_470_), .F2(nn4010), .F3(\coefcal1_divide_inst1_u115_XORCI_1|SUM_net ) );
      defparam ii4114.CONFIG_DATA = 16'hA695;
      defparam ii4114.PLACE_LOCATION = "NONE";
      defparam ii4114.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4115 ( .DX(nn4115), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn4063), .F2(dummy_abc_2861_), .F3(dummy_abc_2862_) );
      defparam ii4115.CONFIG_DATA = 16'h9999;
      defparam ii4115.PLACE_LOCATION = "NONE";
      defparam ii4115.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4116 ( .DX(nn4116), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn4065), .F2(dummy_abc_2863_), .F3(dummy_abc_2864_) );
      defparam ii4116.CONFIG_DATA = 16'h9999;
      defparam ii4116.PLACE_LOCATION = "NONE";
      defparam ii4116.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4117 ( .DX(nn4117), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn4067), .F2(dummy_abc_2865_), .F3(dummy_abc_2866_) );
      defparam ii4117.CONFIG_DATA = 16'h9999;
      defparam ii4117.PLACE_LOCATION = "NONE";
      defparam ii4117.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4118 ( .DX(nn4118), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn4069), .F2(dummy_abc_2867_), .F3(dummy_abc_2868_) );
      defparam ii4118.CONFIG_DATA = 16'h9999;
      defparam ii4118.PLACE_LOCATION = "NONE";
      defparam ii4118.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4119 ( .DX(nn4119), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn4071), .F2(dummy_abc_2869_), .F3(dummy_abc_2870_) );
      defparam ii4119.CONFIG_DATA = 16'h9999;
      defparam ii4119.PLACE_LOCATION = "NONE";
      defparam ii4119.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4120 ( .DX(nn4120), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn4073), .F2(dummy_abc_2871_), .F3(dummy_abc_2872_) );
      defparam ii4120.CONFIG_DATA = 16'h9999;
      defparam ii4120.PLACE_LOCATION = "NONE";
      defparam ii4120.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4121 ( .DX(nn4121), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn4075), .F2(dummy_abc_2873_), .F3(dummy_abc_2874_) );
      defparam ii4121.CONFIG_DATA = 16'h9999;
      defparam ii4121.PLACE_LOCATION = "NONE";
      defparam ii4121.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4122 ( .DX(nn4122), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn4077), .F2(dummy_abc_2875_), .F3(dummy_abc_2876_) );
      defparam ii4122.CONFIG_DATA = 16'h9999;
      defparam ii4122.PLACE_LOCATION = "NONE";
      defparam ii4122.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4123 ( .DX(nn4123), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn4079), .F2(dummy_abc_2877_), .F3(dummy_abc_2878_) );
      defparam ii4123.CONFIG_DATA = 16'h9999;
      defparam ii4123.PLACE_LOCATION = "NONE";
      defparam ii4123.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4124 ( .DX(nn4124), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn4081), .F2(dummy_abc_2879_), .F3(dummy_abc_2880_) );
      defparam ii4124.CONFIG_DATA = 16'h9999;
      defparam ii4124.PLACE_LOCATION = "NONE";
      defparam ii4124.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4125 ( .DX(nn4125), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn4083), .F2(dummy_abc_2881_), .F3(dummy_abc_2882_) );
      defparam ii4125.CONFIG_DATA = 16'h9999;
      defparam ii4125.PLACE_LOCATION = "NONE";
      defparam ii4125.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4126 ( .DX(nn4126), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn4085), .F2(dummy_abc_2883_), .F3(dummy_abc_2884_) );
      defparam ii4126.CONFIG_DATA = 16'h9999;
      defparam ii4126.PLACE_LOCATION = "NONE";
      defparam ii4126.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4127 ( .DX(nn4127), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn4059), .F2(dummy_abc_2885_), .F3(dummy_abc_2886_) );
      defparam ii4127.CONFIG_DATA = 16'h9999;
      defparam ii4127.PLACE_LOCATION = "NONE";
      defparam ii4127.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4128 ( .DX(nn4128), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(dummy_abc_2887_), .F2(dummy_abc_2888_), .F3(dummy_abc_2889_) );
      defparam ii4128.CONFIG_DATA = 16'h5555;
      defparam ii4128.PLACE_LOCATION = "NONE";
      defparam ii4128.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_228_ ( 
        .CA( {a_acc_en_cal1_u137_mac, nn4059, nn4085, nn4083, nn4081, nn4079, 
              nn4077, nn4075, nn4073, nn4071, nn4069, nn4067, nn4065, nn4063, 
              nn4111, nn4110, \coefcal1_xDividend__reg[1]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_169_ ), 
        .DX( {nn4128, nn4127, nn4126, nn4125, nn4124, nn4123, nn4122, nn4121, 
              nn4120, nn4119, nn4118, nn4117, nn4116, nn4115, nn4114, nn4113, 
              nn4112} ), 
        .SUM( {dummy_170_, \coefcal1_divide_inst1_u116_XORCI_15|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_14|SUM_net , \coefcal1_divide_inst1_u116_XORCI_13|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_12|SUM_net , \coefcal1_divide_inst1_u116_XORCI_11|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_10|SUM_net , \coefcal1_divide_inst1_u116_XORCI_9|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_8|SUM_net , \coefcal1_divide_inst1_u116_XORCI_7|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_6|SUM_net , \coefcal1_divide_inst1_u116_XORCI_5|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_4|SUM_net , \coefcal1_divide_inst1_u116_XORCI_3|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_2|SUM_net , \coefcal1_divide_inst1_u116_XORCI_1|SUM_net , 
              \coefcal1_divide_inst1_u116_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4148 ( .DX(nn4148), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(nn4059), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_15|SUM_net ) );
      defparam ii4148.CONFIG_DATA = 16'h202A;
      defparam ii4148.PLACE_LOCATION = "NONE";
      defparam ii4148.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4149 ( .DX(nn4149), .F0(\coefcal1_xDividend__reg[16]|Q_net ), .F1(\coefcal1_xDivisor__reg[16]|Q_net ), .F2(nn4148), .F3(dummy_abc_2890_) );
      defparam ii4149.CONFIG_DATA = 16'h0D0D;
      defparam ii4149.PLACE_LOCATION = "NONE";
      defparam ii4149.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4150 ( .DX(nn4150), .F0(dummy_abc_2891_), .F1(dummy_abc_2892_), .F2(dummy_abc_2893_), .F3(dummy_abc_2894_) );
      defparam ii4150.CONFIG_DATA = 16'hFFFF;
      defparam ii4150.PLACE_LOCATION = "NONE";
      defparam ii4150.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18 ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDividend__reg[16]|Q_net , 
              \coefcal1_xDividend__reg[15]|Q_net , \coefcal1_xDividend__reg[14]|Q_net , 
              \coefcal1_xDividend__reg[13]|Q_net , \coefcal1_xDividend__reg[12]|Q_net , 
              \coefcal1_xDividend__reg[11]|Q_net , \coefcal1_xDividend__reg[10]|Q_net , 
              \coefcal1_xDividend__reg[9]|Q_net , \coefcal1_xDividend__reg[8]|Q_net , 
              \coefcal1_xDividend__reg[7]|Q_net , \coefcal1_xDividend__reg[6]|Q_net , 
              \coefcal1_xDividend__reg[5]|Q_net , \coefcal1_xDividend__reg[4]|Q_net , 
              \coefcal1_xDividend__reg[3]|Q_net , \coefcal1_xDividend__reg[2]|Q_net , 
              \coefcal1_xDividend__reg[1]|Q_net , \coefcal1_xDividend__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_204_ ), 
        .DX( {nn4150, nn4149, nn2918, nn2917, nn2916, nn2915, nn2914, nn2913, 
              nn2912, nn2911, nn2910, nn2909, nn2908, nn2907, nn2906, nn2905, 
              nn2904, nn2903} ), 
        .SUM( {\coefcal1_divide_inst1_u118_XORCI_17|SUM_net , dummy_205_, 
              dummy_206_, dummy_207_, dummy_208_, dummy_209_, dummy_210_, dummy_211_, 
              dummy_212_, dummy_213_, dummy_214_, dummy_215_, dummy_216_, dummy_217_, 
              dummy_218_, dummy_219_, dummy_220_, dummy_221_} )
      );
    CS_LUT4_PRIM ii4171 ( .DX(nn4171), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(\coefcal1_xDivisor__reg[7]|Q_net ), .F2(\coefcal1_xDivisor__reg[8]|Q_net ), .F3(\coefcal1_xDivisor__reg[9]|Q_net ) );
      defparam ii4171.CONFIG_DATA = 16'h0001;
      defparam ii4171.PLACE_LOCATION = "NONE";
      defparam ii4171.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4172 ( .DX(nn4172), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(\coefcal1_xDivisor__reg[2]|Q_net ), .F2(\coefcal1_xDivisor__reg[5]|Q_net ), .F3(nn4171) );
      defparam ii4172.CONFIG_DATA = 16'h0100;
      defparam ii4172.PLACE_LOCATION = "NONE";
      defparam ii4172.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4173 ( .DX(nn4173), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(\coefcal1_xDivisor__reg[15]|Q_net ), .F2(\coefcal1_xDivisor__reg[16]|Q_net ), .F3(\coefcal1_xDivisor__reg[1]|Q_net ) );
      defparam ii4173.CONFIG_DATA = 16'h0001;
      defparam ii4173.PLACE_LOCATION = "NONE";
      defparam ii4173.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4174 ( .DX(nn4174), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(\coefcal1_xDivisor__reg[11]|Q_net ), .F2(\coefcal1_xDivisor__reg[12]|Q_net ), .F3(nn4173) );
      defparam ii4174.CONFIG_DATA = 16'h0100;
      defparam ii4174.PLACE_LOCATION = "NONE";
      defparam ii4174.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4175 ( .DX(nn4175), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(\coefcal1_xDivisor__reg[4]|Q_net ), .F2(nn4172), .F3(nn4174) );
      defparam ii4175.CONFIG_DATA = 16'h1000;
      defparam ii4175.PLACE_LOCATION = "NONE";
      defparam ii4175.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4176 ( .DX(nn4176), .F0(\coefcal1_xDivisor__reg[0]|Q_net ), .F1(nn4175), .F2(dummy_abc_2895_), .F3(dummy_abc_2896_) );
      defparam ii4176.CONFIG_DATA = 16'h4444;
      defparam ii4176.PLACE_LOCATION = "NONE";
      defparam ii4176.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4177 ( .DX(nn4177), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(dummy_abc_2897_), .F3(dummy_abc_2898_) );
      defparam ii4177.CONFIG_DATA = 16'h9999;
      defparam ii4177.PLACE_LOCATION = "NONE";
      defparam ii4177.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4178 ( .DX(nn4178), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(\coefcal1_xDivisor__reg[0]|Q_net ), .F2(\coefcal1_xDivisor__reg[1]|Q_net ), .F3(dummy_489_) );
      defparam ii4178.CONFIG_DATA = 16'hA569;
      defparam ii4178.PLACE_LOCATION = "NONE";
      defparam ii4178.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4179 ( .DX(nn4179), .F0(\coefcal1_xDivisor__reg[2]|Q_net ), .F1(dummy_489_), .F2(nn4110), .F3(\coefcal1_divide_inst1_u116_XORCI_1|SUM_net ) );
      defparam ii4179.CONFIG_DATA = 16'hA695;
      defparam ii4179.PLACE_LOCATION = "NONE";
      defparam ii4179.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4180 ( .DX(nn4180), .F0(\coefcal1_xDivisor__reg[3]|Q_net ), .F1(nn4111), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_2|SUM_net ) );
      defparam ii4180.CONFIG_DATA = 16'h9A95;
      defparam ii4180.PLACE_LOCATION = "NONE";
      defparam ii4180.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4181 ( .DX(nn4181), .F0(\coefcal1_xDivisor__reg[4]|Q_net ), .F1(nn4063), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_3|SUM_net ) );
      defparam ii4181.CONFIG_DATA = 16'h9A95;
      defparam ii4181.PLACE_LOCATION = "NONE";
      defparam ii4181.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4182 ( .DX(nn4182), .F0(\coefcal1_xDivisor__reg[5]|Q_net ), .F1(nn4065), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_4|SUM_net ) );
      defparam ii4182.CONFIG_DATA = 16'h9A95;
      defparam ii4182.PLACE_LOCATION = "NONE";
      defparam ii4182.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4183 ( .DX(nn4183), .F0(\coefcal1_xDivisor__reg[6]|Q_net ), .F1(nn4067), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_5|SUM_net ) );
      defparam ii4183.CONFIG_DATA = 16'h9A95;
      defparam ii4183.PLACE_LOCATION = "NONE";
      defparam ii4183.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4184 ( .DX(nn4184), .F0(\coefcal1_xDivisor__reg[7]|Q_net ), .F1(nn4069), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_6|SUM_net ) );
      defparam ii4184.CONFIG_DATA = 16'h9A95;
      defparam ii4184.PLACE_LOCATION = "NONE";
      defparam ii4184.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4185 ( .DX(nn4185), .F0(\coefcal1_xDivisor__reg[8]|Q_net ), .F1(nn4071), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_7|SUM_net ) );
      defparam ii4185.CONFIG_DATA = 16'h9A95;
      defparam ii4185.PLACE_LOCATION = "NONE";
      defparam ii4185.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4186 ( .DX(nn4186), .F0(\coefcal1_xDivisor__reg[9]|Q_net ), .F1(nn4073), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_8|SUM_net ) );
      defparam ii4186.CONFIG_DATA = 16'h9A95;
      defparam ii4186.PLACE_LOCATION = "NONE";
      defparam ii4186.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4187 ( .DX(nn4187), .F0(\coefcal1_xDivisor__reg[10]|Q_net ), .F1(nn4075), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_9|SUM_net ) );
      defparam ii4187.CONFIG_DATA = 16'h9A95;
      defparam ii4187.PLACE_LOCATION = "NONE";
      defparam ii4187.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4188 ( .DX(nn4188), .F0(\coefcal1_xDivisor__reg[11]|Q_net ), .F1(nn4077), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_10|SUM_net ) );
      defparam ii4188.CONFIG_DATA = 16'h9A95;
      defparam ii4188.PLACE_LOCATION = "NONE";
      defparam ii4188.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4189 ( .DX(nn4189), .F0(\coefcal1_xDivisor__reg[12]|Q_net ), .F1(nn4079), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_11|SUM_net ) );
      defparam ii4189.CONFIG_DATA = 16'h9A95;
      defparam ii4189.PLACE_LOCATION = "NONE";
      defparam ii4189.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4190 ( .DX(nn4190), .F0(\coefcal1_xDivisor__reg[13]|Q_net ), .F1(nn4081), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_12|SUM_net ) );
      defparam ii4190.CONFIG_DATA = 16'h9A95;
      defparam ii4190.PLACE_LOCATION = "NONE";
      defparam ii4190.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4191 ( .DX(nn4191), .F0(\coefcal1_xDivisor__reg[14]|Q_net ), .F1(nn4083), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_13|SUM_net ) );
      defparam ii4191.CONFIG_DATA = 16'h9A95;
      defparam ii4191.PLACE_LOCATION = "NONE";
      defparam ii4191.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4192 ( .DX(nn4192), .F0(\coefcal1_xDivisor__reg[15]|Q_net ), .F1(nn4085), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_14|SUM_net ) );
      defparam ii4192.CONFIG_DATA = 16'h9A95;
      defparam ii4192.PLACE_LOCATION = "NONE";
      defparam ii4192.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4193 ( .DX(nn4193), .F0(\coefcal1_xDivisor__reg[16]|Q_net ), .F1(nn4059), .F2(dummy_489_), .F3(\coefcal1_divide_inst1_u116_XORCI_15|SUM_net ) );
      defparam ii4193.CONFIG_DATA = 16'h9A95;
      defparam ii4193.PLACE_LOCATION = "NONE";
      defparam ii4193.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4194 ( .DX(nn4194), .F0(dummy_abc_2899_), .F1(dummy_abc_2900_), .F2(dummy_abc_2901_), .F3(dummy_abc_2902_) );
      defparam ii4194.CONFIG_DATA = 16'hFFFF;
      defparam ii4194.PLACE_LOCATION = "NONE";
      defparam ii4194.PCK_LOCATION = "NONE";
    scaler_ipc_adder_18 carry_18_244_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \coefcal1_xDivisor__reg[16]|Q_net , 
              \coefcal1_xDivisor__reg[15]|Q_net , \coefcal1_xDivisor__reg[14]|Q_net , 
              \coefcal1_xDivisor__reg[13]|Q_net , \coefcal1_xDivisor__reg[12]|Q_net , 
              \coefcal1_xDivisor__reg[11]|Q_net , \coefcal1_xDivisor__reg[10]|Q_net , 
              \coefcal1_xDivisor__reg[9]|Q_net , \coefcal1_xDivisor__reg[8]|Q_net , 
              \coefcal1_xDivisor__reg[7]|Q_net , \coefcal1_xDivisor__reg[6]|Q_net , 
              \coefcal1_xDivisor__reg[5]|Q_net , \coefcal1_xDivisor__reg[4]|Q_net , 
              \coefcal1_xDivisor__reg[3]|Q_net , \coefcal1_xDivisor__reg[2]|Q_net , 
              \coefcal1_xDivisor__reg[1]|Q_net , \coefcal1_xDivisor__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_508_ ), 
        .DX( {nn4194, nn4193, nn4192, nn4191, nn4190, nn4189, nn4188, nn4187, 
              nn4186, nn4185, nn4184, nn4183, nn4182, nn4181, nn4180, nn4179, 
              nn4178, nn4177} ), 
        .SUM( {\coefcal1_divide_inst1_u150_XORCI_17|SUM_net , dummy_509_, 
              dummy_510_, dummy_511_, dummy_512_, dummy_513_, dummy_514_, dummy_515_, 
              dummy_516_, dummy_517_, dummy_518_, dummy_519_, dummy_520_, dummy_521_, 
              dummy_522_, dummy_523_, dummy_524_, dummy_525_} )
      );
    CS_LUT4_PRIM ii4215 ( .DX(nn4215), .F0(\coefcal1_xDividend__reg[0]|Q_net ), .F1(dummy_508_), .F2(nn4175), .F3(dummy_abc_2903_) );
      defparam ii4215.CONFIG_DATA = 16'h5C5C;
      defparam ii4215.PLACE_LOCATION = "NONE";
      defparam ii4215.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4216 ( .DX(nn4216), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4215) );
      defparam ii4216.CONFIG_DATA = 16'hFFFB;
      defparam ii4216.PLACE_LOCATION = "NONE";
      defparam ii4216.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4217 ( .DX(nn4217), .F0(\cal1_u__reg[0]|Q_net ), .F1(nn4216), .F2(dummy_abc_2904_), .F3(dummy_abc_2905_) );
      defparam ii4217.CONFIG_DATA = 16'h6666;
      defparam ii4217.PLACE_LOCATION = "NONE";
      defparam ii4217.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4218 ( .DX(nn4218), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4215) );
      defparam ii4218.CONFIG_DATA = 16'hFFFB;
      defparam ii4218.PLACE_LOCATION = "NONE";
      defparam ii4218.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4219 ( .DX(nn4219), .F0(\coefcal1_xDividend__reg[1]|Q_net ), .F1(dummy_489_), .F2(nn4175), .F3(dummy_abc_2906_) );
      defparam ii4219.CONFIG_DATA = 16'h5C5C;
      defparam ii4219.PLACE_LOCATION = "NONE";
      defparam ii4219.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4220 ( .DX(nn4220), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4219) );
      defparam ii4220.CONFIG_DATA = 16'h0004;
      defparam ii4220.PLACE_LOCATION = "NONE";
      defparam ii4220.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4221 ( .DX(nn4221), .F0(\coefcal1_xDividend__reg[2]|Q_net ), .F1(dummy_470_), .F2(nn4175), .F3(dummy_abc_2907_) );
      defparam ii4221.CONFIG_DATA = 16'h5C5C;
      defparam ii4221.PLACE_LOCATION = "NONE";
      defparam ii4221.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4222 ( .DX(nn4222), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4221) );
      defparam ii4222.CONFIG_DATA = 16'h0004;
      defparam ii4222.PLACE_LOCATION = "NONE";
      defparam ii4222.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4223 ( .DX(nn4223), .F0(\coefcal1_xDividend__reg[3]|Q_net ), .F1(dummy_451_), .F2(nn4175), .F3(dummy_abc_2908_) );
      defparam ii4223.CONFIG_DATA = 16'h5C5C;
      defparam ii4223.PLACE_LOCATION = "NONE";
      defparam ii4223.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4224 ( .DX(nn4224), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4223) );
      defparam ii4224.CONFIG_DATA = 16'h0004;
      defparam ii4224.PLACE_LOCATION = "NONE";
      defparam ii4224.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4225 ( .DX(nn4225), .F0(\coefcal1_xDividend__reg[4]|Q_net ), .F1(dummy_432_), .F2(nn4175), .F3(dummy_abc_2909_) );
      defparam ii4225.CONFIG_DATA = 16'h5C5C;
      defparam ii4225.PLACE_LOCATION = "NONE";
      defparam ii4225.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4226 ( .DX(nn4226), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4225) );
      defparam ii4226.CONFIG_DATA = 16'h0004;
      defparam ii4226.PLACE_LOCATION = "NONE";
      defparam ii4226.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4227 ( .DX(nn4227), .F0(\coefcal1_xDividend__reg[5]|Q_net ), .F1(dummy_413_), .F2(nn4175), .F3(dummy_abc_2910_) );
      defparam ii4227.CONFIG_DATA = 16'h5C5C;
      defparam ii4227.PLACE_LOCATION = "NONE";
      defparam ii4227.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4228 ( .DX(nn4228), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4227) );
      defparam ii4228.CONFIG_DATA = 16'h0004;
      defparam ii4228.PLACE_LOCATION = "NONE";
      defparam ii4228.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4229 ( .DX(nn4229), .F0(\coefcal1_xDividend__reg[6]|Q_net ), .F1(dummy_394_), .F2(nn4175), .F3(dummy_abc_2911_) );
      defparam ii4229.CONFIG_DATA = 16'h5C5C;
      defparam ii4229.PLACE_LOCATION = "NONE";
      defparam ii4229.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4230 ( .DX(nn4230), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4229) );
      defparam ii4230.CONFIG_DATA = 16'h0004;
      defparam ii4230.PLACE_LOCATION = "NONE";
      defparam ii4230.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4231 ( .DX(nn4231), .F0(\coefcal1_xDividend__reg[7]|Q_net ), .F1(dummy_375_), .F2(nn4175), .F3(dummy_abc_2912_) );
      defparam ii4231.CONFIG_DATA = 16'h5C5C;
      defparam ii4231.PLACE_LOCATION = "NONE";
      defparam ii4231.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4232 ( .DX(nn4232), .F0(rst), .F1(dummy_204_), .F2(nn4176), .F3(nn4231) );
      defparam ii4232.CONFIG_DATA = 16'h0004;
      defparam ii4232.PLACE_LOCATION = "NONE";
      defparam ii4232.PCK_LOCATION = "NONE";
    scaler_ipc_adder_8 carry_8 ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_dinxy_cen_cal1_u137_mac} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_887_ ), 
        .DX( {nn4232, nn4230, nn4228, nn4226, nn4224, nn4222, nn4220, nn4218} ), 
        .SUM( {\coefcal1_u61_XORCI_7|SUM_net , \coefcal1_u61_XORCI_6|SUM_net , 
              \coefcal1_u61_XORCI_5|SUM_net , \coefcal1_u61_XORCI_4|SUM_net , 
              \coefcal1_u61_XORCI_3|SUM_net , \coefcal1_u61_XORCI_2|SUM_net , 
              \coefcal1_u61_XORCI_1|SUM_net , \coefcal1_u61_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4243 ( .DX(nn4243), .F0(\cal1_u__reg[1]|Q_net ), .F1(\coefcal1_u61_XORCI_1|SUM_net ), .F2(dummy_abc_2913_), .F3(dummy_abc_2914_) );
      defparam ii4243.CONFIG_DATA = 16'h6666;
      defparam ii4243.PLACE_LOCATION = "NONE";
      defparam ii4243.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4244 ( .DX(nn4244), .F0(\cal1_u__reg[2]|Q_net ), .F1(\coefcal1_u61_XORCI_2|SUM_net ), .F2(dummy_abc_2915_), .F3(dummy_abc_2916_) );
      defparam ii4244.CONFIG_DATA = 16'h6666;
      defparam ii4244.PLACE_LOCATION = "NONE";
      defparam ii4244.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4245 ( .DX(nn4245), .F0(\cal1_u__reg[3]|Q_net ), .F1(\coefcal1_u61_XORCI_3|SUM_net ), .F2(dummy_abc_2917_), .F3(dummy_abc_2918_) );
      defparam ii4245.CONFIG_DATA = 16'h6666;
      defparam ii4245.PLACE_LOCATION = "NONE";
      defparam ii4245.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4246 ( .DX(nn4246), .F0(\cal1_u__reg[4]|Q_net ), .F1(\coefcal1_u61_XORCI_4|SUM_net ), .F2(dummy_abc_2919_), .F3(dummy_abc_2920_) );
      defparam ii4246.CONFIG_DATA = 16'h6666;
      defparam ii4246.PLACE_LOCATION = "NONE";
      defparam ii4246.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4247 ( .DX(nn4247), .F0(\cal1_u__reg[5]|Q_net ), .F1(\coefcal1_u61_XORCI_5|SUM_net ), .F2(dummy_abc_2921_), .F3(dummy_abc_2922_) );
      defparam ii4247.CONFIG_DATA = 16'h6666;
      defparam ii4247.PLACE_LOCATION = "NONE";
      defparam ii4247.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4248 ( .DX(nn4248), .F0(\cal1_u__reg[6]|Q_net ), .F1(\coefcal1_u61_XORCI_6|SUM_net ), .F2(dummy_abc_2923_), .F3(dummy_abc_2924_) );
      defparam ii4248.CONFIG_DATA = 16'h6666;
      defparam ii4248.PLACE_LOCATION = "NONE";
      defparam ii4248.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4249 ( .DX(nn4249), .F0(\cal1_u__reg[7]|Q_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_abc_2925_), .F3(dummy_abc_2926_) );
      defparam ii4249.CONFIG_DATA = 16'h6666;
      defparam ii4249.PLACE_LOCATION = "NONE";
      defparam ii4249.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4250 ( .DX(nn4250), .F0(\cal1_u__reg[8]|Q_net ), .F1(dummy_abc_2927_), .F2(dummy_abc_2928_), .F3(dummy_abc_2929_) );
      defparam ii4250.CONFIG_DATA = 16'hAAAA;
      defparam ii4250.PLACE_LOCATION = "NONE";
      defparam ii4250.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4251 ( .DX(nn4251), .F0(\cal1_u__reg[9]|Q_net ), .F1(dummy_abc_2930_), .F2(dummy_abc_2931_), .F3(dummy_abc_2932_) );
      defparam ii4251.CONFIG_DATA = 16'hAAAA;
      defparam ii4251.PLACE_LOCATION = "NONE";
      defparam ii4251.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4252 ( .DX(nn4252), .F0(\cal1_u__reg[10]|Q_net ), .F1(dummy_abc_2933_), .F2(dummy_abc_2934_), .F3(dummy_abc_2935_) );
      defparam ii4252.CONFIG_DATA = 16'hAAAA;
      defparam ii4252.PLACE_LOCATION = "NONE";
      defparam ii4252.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4253 ( .DX(nn4253), .F0(\cal1_u__reg[11]|Q_net ), .F1(dummy_abc_2936_), .F2(dummy_abc_2937_), .F3(dummy_abc_2938_) );
      defparam ii4253.CONFIG_DATA = 16'hAAAA;
      defparam ii4253.PLACE_LOCATION = "NONE";
      defparam ii4253.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4254 ( .DX(nn4254), .F0(\cal1_u__reg[12]|Q_net ), .F1(dummy_abc_2939_), .F2(dummy_abc_2940_), .F3(dummy_abc_2941_) );
      defparam ii4254.CONFIG_DATA = 16'hAAAA;
      defparam ii4254.PLACE_LOCATION = "NONE";
      defparam ii4254.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4255 ( .DX(nn4255), .F0(\cal1_u__reg[13]|Q_net ), .F1(dummy_abc_2942_), .F2(dummy_abc_2943_), .F3(dummy_abc_2944_) );
      defparam ii4255.CONFIG_DATA = 16'hAAAA;
      defparam ii4255.PLACE_LOCATION = "NONE";
      defparam ii4255.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4256 ( .DX(nn4256), .F0(\cal1_u__reg[14]|Q_net ), .F1(dummy_abc_2945_), .F2(dummy_abc_2946_), .F3(dummy_abc_2947_) );
      defparam ii4256.CONFIG_DATA = 16'hAAAA;
      defparam ii4256.PLACE_LOCATION = "NONE";
      defparam ii4256.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4257 ( .DX(nn4257), .F0(\cal1_u__reg[15]|Q_net ), .F1(dummy_abc_2948_), .F2(dummy_abc_2949_), .F3(dummy_abc_2950_) );
      defparam ii4257.CONFIG_DATA = 16'hAAAA;
      defparam ii4257.PLACE_LOCATION = "NONE";
      defparam ii4257.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4258 ( .DX(nn4258), .F0(\cal1_u__reg[16]|Q_net ), .F1(dummy_abc_2951_), .F2(dummy_abc_2952_), .F3(dummy_abc_2953_) );
      defparam ii4258.CONFIG_DATA = 16'hAAAA;
      defparam ii4258.PLACE_LOCATION = "NONE";
      defparam ii4258.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17 ( 
        .CA( {\cal1_u__reg[16]|Q_net , \cal1_u__reg[15]|Q_net , 
              \cal1_u__reg[14]|Q_net , \cal1_u__reg[13]|Q_net , \cal1_u__reg[12]|Q_net , 
              \cal1_u__reg[11]|Q_net , \cal1_u__reg[10]|Q_net , \cal1_u__reg[9]|Q_net , 
              \cal1_u__reg[8]|Q_net , \cal1_u__reg[7]|Q_net , \cal1_u__reg[6]|Q_net , 
              \cal1_u__reg[5]|Q_net , \cal1_u__reg[4]|Q_net , \cal1_u__reg[3]|Q_net , 
              \cal1_u__reg[2]|Q_net , \cal1_u__reg[1]|Q_net , \cal1_u__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_139_ ), 
        .DX( {nn4258, nn4257, nn4256, nn4255, nn4254, nn4253, nn4252, nn4251, 
              nn4250, nn4249, nn4248, nn4247, nn4246, nn4245, nn4244, nn4243, 
              nn4217} ), 
        .SUM( {\cal1_u127_XORCI_16|SUM_net , \cal1_u127_XORCI_15|SUM_net , 
              \cal1_u127_XORCI_14|SUM_net , \cal1_u127_XORCI_13|SUM_net , \cal1_u127_XORCI_12|SUM_net , 
              \cal1_u127_XORCI_11|SUM_net , \cal1_u127_XORCI_10|SUM_net , \cal1_u127_XORCI_9|SUM_net , 
              \cal1_u127_XORCI_8|SUM_net , \cal1_u127_XORCI_7|SUM_net , \cal1_u127_XORCI_6|SUM_net , 
              \cal1_u127_XORCI_5|SUM_net , \cal1_u127_XORCI_4|SUM_net , \cal1_u127_XORCI_3|SUM_net , 
              \cal1_u127_XORCI_2|SUM_net , \cal1_u127_XORCI_1|SUM_net , \cal1_u127_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4278 ( .DX(nn4278), .F0(\cal1_u__reg[6]|Q_net ), .F1(\cal1_u__reg[7]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(\cal1_u127_XORCI_7|SUM_net ) );
      defparam ii4278.CONFIG_DATA = 16'h39C6;
      defparam ii4278.PLACE_LOCATION = "NONE";
      defparam ii4278.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4279 ( .DX(nn4279), .F0(\cal1_u__reg[6]|Q_net ), .F1(\cal1_u__reg[7]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(\cal1_u127_XORCI_7|SUM_net ) );
      defparam ii4279.CONFIG_DATA = 16'h08CE;
      defparam ii4279.PLACE_LOCATION = "NONE";
      defparam ii4279.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4280 ( .DX(nn4280), .F0(\cal1_u__reg[8]|Q_net ), .F1(\cal1_u127_XORCI_8|SUM_net ), .F2(nn4278), .F3(nn4279) );
      defparam ii4280.CONFIG_DATA = 16'h0609;
      defparam ii4280.PLACE_LOCATION = "NONE";
      defparam ii4280.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4281 ( .DX(nn4281), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\cal1_u__reg[6]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(nn4280) );
      defparam ii4281.CONFIG_DATA = 16'h96AA;
      defparam ii4281.PLACE_LOCATION = "NONE";
      defparam ii4281.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4282 ( .DX(nn4282), .F0(dummy_36_), .F1(dummy_23_), .F2(nn4281), .F3(dummy_abc_2954_) );
      defparam ii4282.CONFIG_DATA = 16'h8080;
      defparam ii4282.PLACE_LOCATION = "NONE";
      defparam ii4282.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4283 ( .DX(nn4283), .F0(dummy_36_), .F1(dummy_23_), .F2(nn1499), .F3(dummy_abc_2955_) );
      defparam ii4283.CONFIG_DATA = 16'hF7F7;
      defparam ii4283.PLACE_LOCATION = "NONE";
      defparam ii4283.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4284 ( .DX(nn4284), .F0(dummy_49_), .F1(nn1518), .F2(nn4283), .F3(dummy_abc_2956_) );
      defparam ii4284.CONFIG_DATA = 16'hD0D0;
      defparam ii4284.PLACE_LOCATION = "NONE";
      defparam ii4284.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4285 ( .DX(nn4285), .F0(\cal1_ramRdAddr__reg[0]|Q_net ), .F1(\cal1_u__reg[6]|Q_net ), .F2(\cal1_u127_XORCI_6|SUM_net ), .F3(nn4280) );
      defparam ii4285.CONFIG_DATA = 16'h96AA;
      defparam ii4285.PLACE_LOCATION = "NONE";
      defparam ii4285.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4286 ( .DX(nn4286), .F0(\cal1_ramRdAddr__reg[1]|Q_net ), .F1(nn4280), .F2(dummy_abc_2957_), .F3(dummy_abc_2958_) );
      defparam ii4286.CONFIG_DATA = 16'h9999;
      defparam ii4286.PLACE_LOCATION = "NONE";
      defparam ii4286.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4287 ( .DX(nn4287), .F0(\cal1_ramRdAddr__reg[2]|Q_net ), .F1(dummy_abc_2959_), .F2(dummy_abc_2960_), .F3(dummy_abc_2961_) );
      defparam ii4287.CONFIG_DATA = 16'hAAAA;
      defparam ii4287.PLACE_LOCATION = "NONE";
      defparam ii4287.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4288 ( .DX(nn4288), .F0(\cal1_ramRdAddr__reg[3]|Q_net ), .F1(dummy_abc_2962_), .F2(dummy_abc_2963_), .F3(dummy_abc_2964_) );
      defparam ii4288.CONFIG_DATA = 16'hAAAA;
      defparam ii4288.PLACE_LOCATION = "NONE";
      defparam ii4288.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4289 ( .DX(nn4289), .F0(\cal1_ramRdAddr__reg[4]|Q_net ), .F1(dummy_abc_2965_), .F2(dummy_abc_2966_), .F3(dummy_abc_2967_) );
      defparam ii4289.CONFIG_DATA = 16'hAAAA;
      defparam ii4289.PLACE_LOCATION = "NONE";
      defparam ii4289.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4290 ( .DX(nn4290), .F0(\cal1_ramRdAddr__reg[5]|Q_net ), .F1(dummy_abc_2968_), .F2(dummy_abc_2969_), .F3(dummy_abc_2970_) );
      defparam ii4290.CONFIG_DATA = 16'hAAAA;
      defparam ii4290.PLACE_LOCATION = "NONE";
      defparam ii4290.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4291 ( .DX(nn4291), .F0(\cal1_ramRdAddr__reg[6]|Q_net ), .F1(dummy_abc_2971_), .F2(dummy_abc_2972_), .F3(dummy_abc_2973_) );
      defparam ii4291.CONFIG_DATA = 16'hAAAA;
      defparam ii4291.PLACE_LOCATION = "NONE";
      defparam ii4291.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4292 ( .DX(nn4292), .F0(\cal1_ramRdAddr__reg[7]|Q_net ), .F1(dummy_abc_2974_), .F2(dummy_abc_2975_), .F3(dummy_abc_2976_) );
      defparam ii4292.CONFIG_DATA = 16'hAAAA;
      defparam ii4292.PLACE_LOCATION = "NONE";
      defparam ii4292.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4293 ( .DX(nn4293), .F0(\cal1_ramRdAddr__reg[8]|Q_net ), .F1(dummy_abc_2977_), .F2(dummy_abc_2978_), .F3(dummy_abc_2979_) );
      defparam ii4293.CONFIG_DATA = 16'hAAAA;
      defparam ii4293.PLACE_LOCATION = "NONE";
      defparam ii4293.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4294 ( .DX(nn4294), .F0(\cal1_ramRdAddr__reg[9]|Q_net ), .F1(dummy_abc_2980_), .F2(dummy_abc_2981_), .F3(dummy_abc_2982_) );
      defparam ii4294.CONFIG_DATA = 16'hAAAA;
      defparam ii4294.PLACE_LOCATION = "NONE";
      defparam ii4294.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4295 ( .DX(nn4295), .F0(\cal1_ramRdAddr__reg[10]|Q_net ), .F1(dummy_abc_2983_), .F2(dummy_abc_2984_), .F3(dummy_abc_2985_) );
      defparam ii4295.CONFIG_DATA = 16'hAAAA;
      defparam ii4295.PLACE_LOCATION = "NONE";
      defparam ii4295.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_199_ ( 
        .CA( {\cal1_ramRdAddr__reg[10]|Q_net , \cal1_ramRdAddr__reg[9]|Q_net , 
              \cal1_ramRdAddr__reg[8]|Q_net , \cal1_ramRdAddr__reg[7]|Q_net , 
              \cal1_ramRdAddr__reg[6]|Q_net , \cal1_ramRdAddr__reg[5]|Q_net , 
              \cal1_ramRdAddr__reg[4]|Q_net , \cal1_ramRdAddr__reg[3]|Q_net , 
              \cal1_ramRdAddr__reg[2]|Q_net , \cal1_ramRdAddr__reg[1]|Q_net , 
              \cal1_ramRdAddr__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_14_ ), 
        .DX( {nn4295, nn4294, nn4293, nn4292, nn4291, nn4290, nn4289, nn4288, 
              nn4287, nn4286, nn4285} ), 
        .SUM( {\cal1_u130_XORCI_10|SUM_net , \cal1_u130_XORCI_9|SUM_net , 
              \cal1_u130_XORCI_8|SUM_net , \cal1_u130_XORCI_7|SUM_net , \cal1_u130_XORCI_6|SUM_net , 
              \cal1_u130_XORCI_5|SUM_net , \cal1_u130_XORCI_4|SUM_net , \cal1_u130_XORCI_3|SUM_net , 
              \cal1_u130_XORCI_2|SUM_net , \cal1_u130_XORCI_1|SUM_net , \cal1_u130_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4309 ( .DX(nn4309), .F0(\cal1_u130_XORCI_10|SUM_net ), .F1(nn1518), .F2(dummy_abc_2986_), .F3(dummy_abc_2987_) );
      defparam ii4309.CONFIG_DATA = 16'h2222;
      defparam ii4309.PLACE_LOCATION = "NONE";
      defparam ii4309.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4310 ( .DX(nn4310), .F0(\cal1_u130_XORCI_1|SUM_net ), .F1(nn1518), .F2(dummy_abc_2988_), .F3(dummy_abc_2989_) );
      defparam ii4310.CONFIG_DATA = 16'h2222;
      defparam ii4310.PLACE_LOCATION = "NONE";
      defparam ii4310.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4311 ( .DX(nn4311), .F0(\cal1_u130_XORCI_2|SUM_net ), .F1(nn1518), .F2(dummy_abc_2990_), .F3(dummy_abc_2991_) );
      defparam ii4311.CONFIG_DATA = 16'h2222;
      defparam ii4311.PLACE_LOCATION = "NONE";
      defparam ii4311.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4312 ( .DX(nn4312), .F0(\cal1_u130_XORCI_3|SUM_net ), .F1(nn1518), .F2(dummy_abc_2992_), .F3(dummy_abc_2993_) );
      defparam ii4312.CONFIG_DATA = 16'h2222;
      defparam ii4312.PLACE_LOCATION = "NONE";
      defparam ii4312.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4313 ( .DX(nn4313), .F0(\cal1_u130_XORCI_4|SUM_net ), .F1(nn1518), .F2(dummy_abc_2994_), .F3(dummy_abc_2995_) );
      defparam ii4313.CONFIG_DATA = 16'h2222;
      defparam ii4313.PLACE_LOCATION = "NONE";
      defparam ii4313.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4314 ( .DX(nn4314), .F0(\cal1_u130_XORCI_5|SUM_net ), .F1(nn1518), .F2(dummy_abc_2996_), .F3(dummy_abc_2997_) );
      defparam ii4314.CONFIG_DATA = 16'h2222;
      defparam ii4314.PLACE_LOCATION = "NONE";
      defparam ii4314.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4315 ( .DX(nn4315), .F0(\cal1_u130_XORCI_6|SUM_net ), .F1(nn1518), .F2(dummy_abc_2998_), .F3(dummy_abc_2999_) );
      defparam ii4315.CONFIG_DATA = 16'h2222;
      defparam ii4315.PLACE_LOCATION = "NONE";
      defparam ii4315.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4316 ( .DX(nn4316), .F0(\cal1_u130_XORCI_7|SUM_net ), .F1(nn1518), .F2(dummy_abc_3000_), .F3(dummy_abc_3001_) );
      defparam ii4316.CONFIG_DATA = 16'h2222;
      defparam ii4316.PLACE_LOCATION = "NONE";
      defparam ii4316.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4317 ( .DX(nn4317), .F0(\cal1_u130_XORCI_8|SUM_net ), .F1(nn1518), .F2(dummy_abc_3002_), .F3(dummy_abc_3003_) );
      defparam ii4317.CONFIG_DATA = 16'h2222;
      defparam ii4317.PLACE_LOCATION = "NONE";
      defparam ii4317.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4318 ( .DX(nn4318), .F0(\cal1_u130_XORCI_9|SUM_net ), .F1(nn1518), .F2(dummy_abc_3004_), .F3(dummy_abc_3005_) );
      defparam ii4318.CONFIG_DATA = 16'h2222;
      defparam ii4318.PLACE_LOCATION = "NONE";
      defparam ii4318.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4319 ( .DX(nn4319), .F0(\cal1_u__reg[0]|Q_net ), .F1(nn4216), .F2(dummy_abc_3006_), .F3(dummy_abc_3007_) );
      defparam ii4319.CONFIG_DATA = 16'h6666;
      defparam ii4319.PLACE_LOCATION = "NONE";
      defparam ii4319.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4320 ( .DX(nn4320), .F0(nn4319), .F1(nn1518), .F2(dummy_abc_3008_), .F3(dummy_abc_3009_) );
      defparam ii4320.CONFIG_DATA = 16'h2222;
      defparam ii4320.PLACE_LOCATION = "NONE";
      defparam ii4320.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4321 ( .DX(nn4321), .F0(\cal1_u127_XORCI_10|SUM_net ), .F1(nn1518), .F2(dummy_abc_3010_), .F3(dummy_abc_3011_) );
      defparam ii4321.CONFIG_DATA = 16'h2222;
      defparam ii4321.PLACE_LOCATION = "NONE";
      defparam ii4321.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4322 ( .DX(nn4322), .F0(\cal1_u127_XORCI_11|SUM_net ), .F1(nn1518), .F2(dummy_abc_3012_), .F3(dummy_abc_3013_) );
      defparam ii4322.CONFIG_DATA = 16'h2222;
      defparam ii4322.PLACE_LOCATION = "NONE";
      defparam ii4322.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4323 ( .DX(nn4323), .F0(\cal1_u127_XORCI_12|SUM_net ), .F1(nn1518), .F2(dummy_abc_3014_), .F3(dummy_abc_3015_) );
      defparam ii4323.CONFIG_DATA = 16'h2222;
      defparam ii4323.PLACE_LOCATION = "NONE";
      defparam ii4323.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4324 ( .DX(nn4324), .F0(\cal1_u127_XORCI_13|SUM_net ), .F1(nn1518), .F2(dummy_abc_3016_), .F3(dummy_abc_3017_) );
      defparam ii4324.CONFIG_DATA = 16'h2222;
      defparam ii4324.PLACE_LOCATION = "NONE";
      defparam ii4324.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4325 ( .DX(nn4325), .F0(\cal1_u127_XORCI_14|SUM_net ), .F1(nn1518), .F2(dummy_abc_3018_), .F3(dummy_abc_3019_) );
      defparam ii4325.CONFIG_DATA = 16'h2222;
      defparam ii4325.PLACE_LOCATION = "NONE";
      defparam ii4325.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4326 ( .DX(nn4326), .F0(\cal1_u127_XORCI_15|SUM_net ), .F1(nn1518), .F2(dummy_abc_3020_), .F3(dummy_abc_3021_) );
      defparam ii4326.CONFIG_DATA = 16'h2222;
      defparam ii4326.PLACE_LOCATION = "NONE";
      defparam ii4326.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4327 ( .DX(nn4327), .F0(\cal1_u127_XORCI_16|SUM_net ), .F1(nn1518), .F2(dummy_abc_3022_), .F3(dummy_abc_3023_) );
      defparam ii4327.CONFIG_DATA = 16'h2222;
      defparam ii4327.PLACE_LOCATION = "NONE";
      defparam ii4327.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4328 ( .DX(nn4328), .F0(\cal1_u127_XORCI_1|SUM_net ), .F1(nn1518), .F2(dummy_abc_3024_), .F3(dummy_abc_3025_) );
      defparam ii4328.CONFIG_DATA = 16'h2222;
      defparam ii4328.PLACE_LOCATION = "NONE";
      defparam ii4328.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4329 ( .DX(nn4329), .F0(\cal1_u127_XORCI_2|SUM_net ), .F1(nn1518), .F2(dummy_abc_3026_), .F3(dummy_abc_3027_) );
      defparam ii4329.CONFIG_DATA = 16'h2222;
      defparam ii4329.PLACE_LOCATION = "NONE";
      defparam ii4329.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4330 ( .DX(nn4330), .F0(\cal1_u127_XORCI_3|SUM_net ), .F1(nn1518), .F2(dummy_abc_3028_), .F3(dummy_abc_3029_) );
      defparam ii4330.CONFIG_DATA = 16'h2222;
      defparam ii4330.PLACE_LOCATION = "NONE";
      defparam ii4330.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4331 ( .DX(nn4331), .F0(\cal1_u127_XORCI_4|SUM_net ), .F1(nn1518), .F2(dummy_abc_3030_), .F3(dummy_abc_3031_) );
      defparam ii4331.CONFIG_DATA = 16'h2222;
      defparam ii4331.PLACE_LOCATION = "NONE";
      defparam ii4331.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4332 ( .DX(nn4332), .F0(\cal1_u127_XORCI_5|SUM_net ), .F1(nn1518), .F2(dummy_abc_3032_), .F3(dummy_abc_3033_) );
      defparam ii4332.CONFIG_DATA = 16'h2222;
      defparam ii4332.PLACE_LOCATION = "NONE";
      defparam ii4332.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4333 ( .DX(nn4333), .F0(\cal1_u127_XORCI_6|SUM_net ), .F1(nn1518), .F2(dummy_abc_3034_), .F3(dummy_abc_3035_) );
      defparam ii4333.CONFIG_DATA = 16'h2222;
      defparam ii4333.PLACE_LOCATION = "NONE";
      defparam ii4333.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4334 ( .DX(nn4334), .F0(\cal1_u127_XORCI_7|SUM_net ), .F1(nn1518), .F2(dummy_abc_3036_), .F3(dummy_abc_3037_) );
      defparam ii4334.CONFIG_DATA = 16'h2222;
      defparam ii4334.PLACE_LOCATION = "NONE";
      defparam ii4334.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4335 ( .DX(nn4335), .F0(\cal1_u127_XORCI_8|SUM_net ), .F1(nn1518), .F2(dummy_abc_3038_), .F3(dummy_abc_3039_) );
      defparam ii4335.CONFIG_DATA = 16'h2222;
      defparam ii4335.PLACE_LOCATION = "NONE";
      defparam ii4335.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4336 ( .DX(nn4336), .F0(\cal1_u127_XORCI_9|SUM_net ), .F1(nn1518), .F2(dummy_abc_3040_), .F3(dummy_abc_3041_) );
      defparam ii4336.CONFIG_DATA = 16'h2222;
      defparam ii4336.PLACE_LOCATION = "NONE";
      defparam ii4336.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4337 ( .DX(nn4337), .F0(\cal1_v__reg[0]|Q_net ), .F1(nn2835), .F2(dummy_abc_3042_), .F3(dummy_abc_3043_) );
      defparam ii4337.CONFIG_DATA = 16'h6666;
      defparam ii4337.PLACE_LOCATION = "NONE";
      defparam ii4337.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4338 ( .DX(nn4338), .F0(dummy_36_), .F1(nn4337), .F2(dummy_abc_3044_), .F3(dummy_abc_3045_) );
      defparam ii4338.CONFIG_DATA = 16'h8888;
      defparam ii4338.PLACE_LOCATION = "NONE";
      defparam ii4338.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4339 ( .DX(nn4339), .F0(dummy_36_), .F1(\cal1_u128_XORCI_10|SUM_net ), .F2(dummy_abc_3046_), .F3(dummy_abc_3047_) );
      defparam ii4339.CONFIG_DATA = 16'h8888;
      defparam ii4339.PLACE_LOCATION = "NONE";
      defparam ii4339.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4340 ( .DX(nn4340), .F0(dummy_36_), .F1(\cal1_u128_XORCI_11|SUM_net ), .F2(dummy_abc_3048_), .F3(dummy_abc_3049_) );
      defparam ii4340.CONFIG_DATA = 16'h8888;
      defparam ii4340.PLACE_LOCATION = "NONE";
      defparam ii4340.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4341 ( .DX(nn4341), .F0(dummy_36_), .F1(\cal1_u128_XORCI_12|SUM_net ), .F2(dummy_abc_3050_), .F3(dummy_abc_3051_) );
      defparam ii4341.CONFIG_DATA = 16'h8888;
      defparam ii4341.PLACE_LOCATION = "NONE";
      defparam ii4341.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4342 ( .DX(nn4342), .F0(dummy_36_), .F1(\cal1_u128_XORCI_13|SUM_net ), .F2(dummy_abc_3052_), .F3(dummy_abc_3053_) );
      defparam ii4342.CONFIG_DATA = 16'h8888;
      defparam ii4342.PLACE_LOCATION = "NONE";
      defparam ii4342.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4343 ( .DX(nn4343), .F0(dummy_36_), .F1(\cal1_u128_XORCI_14|SUM_net ), .F2(dummy_abc_3054_), .F3(dummy_abc_3055_) );
      defparam ii4343.CONFIG_DATA = 16'h8888;
      defparam ii4343.PLACE_LOCATION = "NONE";
      defparam ii4343.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4344 ( .DX(nn4344), .F0(dummy_36_), .F1(\cal1_u128_XORCI_15|SUM_net ), .F2(dummy_abc_3056_), .F3(dummy_abc_3057_) );
      defparam ii4344.CONFIG_DATA = 16'h8888;
      defparam ii4344.PLACE_LOCATION = "NONE";
      defparam ii4344.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4345 ( .DX(nn4345), .F0(dummy_36_), .F1(\cal1_u128_XORCI_16|SUM_net ), .F2(dummy_abc_3058_), .F3(dummy_abc_3059_) );
      defparam ii4345.CONFIG_DATA = 16'h8888;
      defparam ii4345.PLACE_LOCATION = "NONE";
      defparam ii4345.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4346 ( .DX(nn4346), .F0(dummy_36_), .F1(\cal1_u128_XORCI_1|SUM_net ), .F2(dummy_abc_3060_), .F3(dummy_abc_3061_) );
      defparam ii4346.CONFIG_DATA = 16'h8888;
      defparam ii4346.PLACE_LOCATION = "NONE";
      defparam ii4346.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4347 ( .DX(nn4347), .F0(dummy_36_), .F1(\cal1_u128_XORCI_2|SUM_net ), .F2(dummy_abc_3062_), .F3(dummy_abc_3063_) );
      defparam ii4347.CONFIG_DATA = 16'h8888;
      defparam ii4347.PLACE_LOCATION = "NONE";
      defparam ii4347.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4348 ( .DX(nn4348), .F0(dummy_36_), .F1(\cal1_u128_XORCI_3|SUM_net ), .F2(dummy_abc_3064_), .F3(dummy_abc_3065_) );
      defparam ii4348.CONFIG_DATA = 16'h8888;
      defparam ii4348.PLACE_LOCATION = "NONE";
      defparam ii4348.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4349 ( .DX(nn4349), .F0(dummy_36_), .F1(\cal1_u128_XORCI_4|SUM_net ), .F2(dummy_abc_3066_), .F3(dummy_abc_3067_) );
      defparam ii4349.CONFIG_DATA = 16'h8888;
      defparam ii4349.PLACE_LOCATION = "NONE";
      defparam ii4349.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4350 ( .DX(nn4350), .F0(dummy_36_), .F1(\cal1_u128_XORCI_5|SUM_net ), .F2(dummy_abc_3068_), .F3(dummy_abc_3069_) );
      defparam ii4350.CONFIG_DATA = 16'h8888;
      defparam ii4350.PLACE_LOCATION = "NONE";
      defparam ii4350.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4351 ( .DX(nn4351), .F0(dummy_36_), .F1(\cal1_u128_XORCI_6|SUM_net ), .F2(dummy_abc_3070_), .F3(dummy_abc_3071_) );
      defparam ii4351.CONFIG_DATA = 16'h8888;
      defparam ii4351.PLACE_LOCATION = "NONE";
      defparam ii4351.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4352 ( .DX(nn4352), .F0(dummy_36_), .F1(\cal1_u128_XORCI_7|SUM_net ), .F2(dummy_abc_3072_), .F3(dummy_abc_3073_) );
      defparam ii4352.CONFIG_DATA = 16'h8888;
      defparam ii4352.PLACE_LOCATION = "NONE";
      defparam ii4352.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4353 ( .DX(nn4353), .F0(dummy_36_), .F1(\cal1_u128_XORCI_8|SUM_net ), .F2(dummy_abc_3074_), .F3(dummy_abc_3075_) );
      defparam ii4353.CONFIG_DATA = 16'h8888;
      defparam ii4353.PLACE_LOCATION = "NONE";
      defparam ii4353.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4354 ( .DX(nn4354), .F0(dummy_36_), .F1(\cal1_u128_XORCI_9|SUM_net ), .F2(dummy_abc_3076_), .F3(dummy_abc_3077_) );
      defparam ii4354.CONFIG_DATA = 16'h8888;
      defparam ii4354.PLACE_LOCATION = "NONE";
      defparam ii4354.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4355 ( .DX(nn4355), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(nn1518), .F2(dummy_abc_3078_), .F3(dummy_abc_3079_) );
      defparam ii4355.CONFIG_DATA = 16'h1111;
      defparam ii4355.PLACE_LOCATION = "NONE";
      defparam ii4355.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4356 ( .DX(nn4356), .F0(\cal1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_3080_), .F2(dummy_abc_3081_), .F3(dummy_abc_3082_) );
      defparam ii4356.CONFIG_DATA = 16'h5555;
      defparam ii4356.PLACE_LOCATION = "NONE";
      defparam ii4356.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4357 ( .DX(nn4357), .F0(\cal1_xAddress__reg[1]|Q_net ), .F1(dummy_abc_3083_), .F2(dummy_abc_3084_), .F3(dummy_abc_3085_) );
      defparam ii4357.CONFIG_DATA = 16'hAAAA;
      defparam ii4357.PLACE_LOCATION = "NONE";
      defparam ii4357.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4358 ( .DX(nn4358), .F0(\cal1_xAddress__reg[2]|Q_net ), .F1(dummy_abc_3086_), .F2(dummy_abc_3087_), .F3(dummy_abc_3088_) );
      defparam ii4358.CONFIG_DATA = 16'hAAAA;
      defparam ii4358.PLACE_LOCATION = "NONE";
      defparam ii4358.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4359 ( .DX(nn4359), .F0(\cal1_xAddress__reg[3]|Q_net ), .F1(dummy_abc_3089_), .F2(dummy_abc_3090_), .F3(dummy_abc_3091_) );
      defparam ii4359.CONFIG_DATA = 16'hAAAA;
      defparam ii4359.PLACE_LOCATION = "NONE";
      defparam ii4359.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4360 ( .DX(nn4360), .F0(\cal1_xAddress__reg[4]|Q_net ), .F1(dummy_abc_3092_), .F2(dummy_abc_3093_), .F3(dummy_abc_3094_) );
      defparam ii4360.CONFIG_DATA = 16'hAAAA;
      defparam ii4360.PLACE_LOCATION = "NONE";
      defparam ii4360.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4361 ( .DX(nn4361), .F0(\cal1_xAddress__reg[5]|Q_net ), .F1(dummy_abc_3095_), .F2(dummy_abc_3096_), .F3(dummy_abc_3097_) );
      defparam ii4361.CONFIG_DATA = 16'hAAAA;
      defparam ii4361.PLACE_LOCATION = "NONE";
      defparam ii4361.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4362 ( .DX(nn4362), .F0(\cal1_xAddress__reg[6]|Q_net ), .F1(dummy_abc_3098_), .F2(dummy_abc_3099_), .F3(dummy_abc_3100_) );
      defparam ii4362.CONFIG_DATA = 16'hAAAA;
      defparam ii4362.PLACE_LOCATION = "NONE";
      defparam ii4362.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4363 ( .DX(nn4363), .F0(\cal1_xAddress__reg[7]|Q_net ), .F1(dummy_abc_3101_), .F2(dummy_abc_3102_), .F3(dummy_abc_3103_) );
      defparam ii4363.CONFIG_DATA = 16'hAAAA;
      defparam ii4363.PLACE_LOCATION = "NONE";
      defparam ii4363.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4364 ( .DX(nn4364), .F0(\cal1_xAddress__reg[8]|Q_net ), .F1(dummy_abc_3104_), .F2(dummy_abc_3105_), .F3(dummy_abc_3106_) );
      defparam ii4364.CONFIG_DATA = 16'hAAAA;
      defparam ii4364.PLACE_LOCATION = "NONE";
      defparam ii4364.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4365 ( .DX(nn4365), .F0(\cal1_xAddress__reg[9]|Q_net ), .F1(dummy_abc_3107_), .F2(dummy_abc_3108_), .F3(dummy_abc_3109_) );
      defparam ii4365.CONFIG_DATA = 16'hAAAA;
      defparam ii4365.PLACE_LOCATION = "NONE";
      defparam ii4365.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4366 ( .DX(nn4366), .F0(\cal1_xAddress__reg[10]|Q_net ), .F1(dummy_abc_3110_), .F2(dummy_abc_3111_), .F3(dummy_abc_3112_) );
      defparam ii4366.CONFIG_DATA = 16'hAAAA;
      defparam ii4366.PLACE_LOCATION = "NONE";
      defparam ii4366.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_200_ ( 
        .CA( {\cal1_xAddress__reg[10]|Q_net , \cal1_xAddress__reg[9]|Q_net , 
              \cal1_xAddress__reg[8]|Q_net , \cal1_xAddress__reg[7]|Q_net , 
              \cal1_xAddress__reg[6]|Q_net , \cal1_xAddress__reg[5]|Q_net , 
              \cal1_xAddress__reg[4]|Q_net , \cal1_xAddress__reg[3]|Q_net , 
              \cal1_xAddress__reg[2]|Q_net , \cal1_xAddress__reg[1]|Q_net , 
              \cal1_xAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_15_ ), 
        .DX( {nn4366, nn4365, nn4364, nn4363, nn4362, nn4361, nn4360, nn4359, 
              nn4358, nn4357, nn4356} ), 
        .SUM( {\cal1_u131_XORCI_10|SUM_net , \cal1_u131_XORCI_9|SUM_net , 
              \cal1_u131_XORCI_8|SUM_net , \cal1_u131_XORCI_7|SUM_net , \cal1_u131_XORCI_6|SUM_net , 
              \cal1_u131_XORCI_5|SUM_net , \cal1_u131_XORCI_4|SUM_net , \cal1_u131_XORCI_3|SUM_net , 
              \cal1_u131_XORCI_2|SUM_net , \cal1_u131_XORCI_1|SUM_net , \cal1_u131_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4380 ( .DX(nn4380), .F0(\cal1_u131_XORCI_10|SUM_net ), .F1(nn1518), .F2(dummy_abc_3113_), .F3(dummy_abc_3114_) );
      defparam ii4380.CONFIG_DATA = 16'h2222;
      defparam ii4380.PLACE_LOCATION = "NONE";
      defparam ii4380.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4381 ( .DX(nn4381), .F0(\cal1_u131_XORCI_1|SUM_net ), .F1(nn1518), .F2(dummy_abc_3115_), .F3(dummy_abc_3116_) );
      defparam ii4381.CONFIG_DATA = 16'h2222;
      defparam ii4381.PLACE_LOCATION = "NONE";
      defparam ii4381.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4382 ( .DX(nn4382), .F0(\cal1_u131_XORCI_2|SUM_net ), .F1(nn1518), .F2(dummy_abc_3117_), .F3(dummy_abc_3118_) );
      defparam ii4382.CONFIG_DATA = 16'h2222;
      defparam ii4382.PLACE_LOCATION = "NONE";
      defparam ii4382.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4383 ( .DX(nn4383), .F0(\cal1_u131_XORCI_3|SUM_net ), .F1(nn1518), .F2(dummy_abc_3119_), .F3(dummy_abc_3120_) );
      defparam ii4383.CONFIG_DATA = 16'h2222;
      defparam ii4383.PLACE_LOCATION = "NONE";
      defparam ii4383.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4384 ( .DX(nn4384), .F0(\cal1_u131_XORCI_4|SUM_net ), .F1(nn1518), .F2(dummy_abc_3121_), .F3(dummy_abc_3122_) );
      defparam ii4384.CONFIG_DATA = 16'h2222;
      defparam ii4384.PLACE_LOCATION = "NONE";
      defparam ii4384.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4385 ( .DX(nn4385), .F0(\cal1_u131_XORCI_5|SUM_net ), .F1(nn1518), .F2(dummy_abc_3123_), .F3(dummy_abc_3124_) );
      defparam ii4385.CONFIG_DATA = 16'h2222;
      defparam ii4385.PLACE_LOCATION = "NONE";
      defparam ii4385.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4386 ( .DX(nn4386), .F0(\cal1_u131_XORCI_6|SUM_net ), .F1(nn1518), .F2(dummy_abc_3125_), .F3(dummy_abc_3126_) );
      defparam ii4386.CONFIG_DATA = 16'h2222;
      defparam ii4386.PLACE_LOCATION = "NONE";
      defparam ii4386.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4387 ( .DX(nn4387), .F0(\cal1_u131_XORCI_7|SUM_net ), .F1(nn1518), .F2(dummy_abc_3127_), .F3(dummy_abc_3128_) );
      defparam ii4387.CONFIG_DATA = 16'h2222;
      defparam ii4387.PLACE_LOCATION = "NONE";
      defparam ii4387.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4388 ( .DX(nn4388), .F0(\cal1_u131_XORCI_8|SUM_net ), .F1(nn1518), .F2(dummy_abc_3129_), .F3(dummy_abc_3130_) );
      defparam ii4388.CONFIG_DATA = 16'h2222;
      defparam ii4388.PLACE_LOCATION = "NONE";
      defparam ii4388.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4389 ( .DX(nn4389), .F0(\cal1_u131_XORCI_9|SUM_net ), .F1(nn1518), .F2(dummy_abc_3131_), .F3(dummy_abc_3132_) );
      defparam ii4389.CONFIG_DATA = 16'h2222;
      defparam ii4389.PLACE_LOCATION = "NONE";
      defparam ii4389.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4390 ( .DX(nn4390), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(dummy_36_), .F2(dummy_abc_3133_), .F3(dummy_abc_3134_) );
      defparam ii4390.CONFIG_DATA = 16'h7777;
      defparam ii4390.PLACE_LOCATION = "NONE";
      defparam ii4390.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4391 ( .DX(nn4391), .F0(\cal1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_3135_), .F2(dummy_abc_3136_), .F3(dummy_abc_3137_) );
      defparam ii4391.CONFIG_DATA = 16'h5555;
      defparam ii4391.PLACE_LOCATION = "NONE";
      defparam ii4391.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4392 ( .DX(nn4392), .F0(\cal1_yAddress__reg[1]|Q_net ), .F1(dummy_abc_3138_), .F2(dummy_abc_3139_), .F3(dummy_abc_3140_) );
      defparam ii4392.CONFIG_DATA = 16'hAAAA;
      defparam ii4392.PLACE_LOCATION = "NONE";
      defparam ii4392.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4393 ( .DX(nn4393), .F0(\cal1_yAddress__reg[2]|Q_net ), .F1(dummy_abc_3141_), .F2(dummy_abc_3142_), .F3(dummy_abc_3143_) );
      defparam ii4393.CONFIG_DATA = 16'hAAAA;
      defparam ii4393.PLACE_LOCATION = "NONE";
      defparam ii4393.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4394 ( .DX(nn4394), .F0(\cal1_yAddress__reg[3]|Q_net ), .F1(dummy_abc_3144_), .F2(dummy_abc_3145_), .F3(dummy_abc_3146_) );
      defparam ii4394.CONFIG_DATA = 16'hAAAA;
      defparam ii4394.PLACE_LOCATION = "NONE";
      defparam ii4394.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4395 ( .DX(nn4395), .F0(\cal1_yAddress__reg[4]|Q_net ), .F1(dummy_abc_3147_), .F2(dummy_abc_3148_), .F3(dummy_abc_3149_) );
      defparam ii4395.CONFIG_DATA = 16'hAAAA;
      defparam ii4395.PLACE_LOCATION = "NONE";
      defparam ii4395.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4396 ( .DX(nn4396), .F0(\cal1_yAddress__reg[5]|Q_net ), .F1(dummy_abc_3150_), .F2(dummy_abc_3151_), .F3(dummy_abc_3152_) );
      defparam ii4396.CONFIG_DATA = 16'hAAAA;
      defparam ii4396.PLACE_LOCATION = "NONE";
      defparam ii4396.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4397 ( .DX(nn4397), .F0(\cal1_yAddress__reg[6]|Q_net ), .F1(dummy_abc_3153_), .F2(dummy_abc_3154_), .F3(dummy_abc_3155_) );
      defparam ii4397.CONFIG_DATA = 16'hAAAA;
      defparam ii4397.PLACE_LOCATION = "NONE";
      defparam ii4397.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4398 ( .DX(nn4398), .F0(\cal1_yAddress__reg[7]|Q_net ), .F1(dummy_abc_3156_), .F2(dummy_abc_3157_), .F3(dummy_abc_3158_) );
      defparam ii4398.CONFIG_DATA = 16'hAAAA;
      defparam ii4398.PLACE_LOCATION = "NONE";
      defparam ii4398.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4399 ( .DX(nn4399), .F0(\cal1_yAddress__reg[8]|Q_net ), .F1(dummy_abc_3159_), .F2(dummy_abc_3160_), .F3(dummy_abc_3161_) );
      defparam ii4399.CONFIG_DATA = 16'hAAAA;
      defparam ii4399.PLACE_LOCATION = "NONE";
      defparam ii4399.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4400 ( .DX(nn4400), .F0(\cal1_yAddress__reg[9]|Q_net ), .F1(dummy_abc_3162_), .F2(dummy_abc_3163_), .F3(dummy_abc_3164_) );
      defparam ii4400.CONFIG_DATA = 16'hAAAA;
      defparam ii4400.PLACE_LOCATION = "NONE";
      defparam ii4400.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4401 ( .DX(nn4401), .F0(\cal1_yAddress__reg[10]|Q_net ), .F1(dummy_abc_3165_), .F2(dummy_abc_3166_), .F3(dummy_abc_3167_) );
      defparam ii4401.CONFIG_DATA = 16'hAAAA;
      defparam ii4401.PLACE_LOCATION = "NONE";
      defparam ii4401.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_201_ ( 
        .CA( {\cal1_yAddress__reg[10]|Q_net , \cal1_yAddress__reg[9]|Q_net , 
              \cal1_yAddress__reg[8]|Q_net , \cal1_yAddress__reg[7]|Q_net , 
              \cal1_yAddress__reg[6]|Q_net , \cal1_yAddress__reg[5]|Q_net , 
              \cal1_yAddress__reg[4]|Q_net , \cal1_yAddress__reg[3]|Q_net , 
              \cal1_yAddress__reg[2]|Q_net , \cal1_yAddress__reg[1]|Q_net , 
              \cal1_yAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_16_ ), 
        .DX( {nn4401, nn4400, nn4399, nn4398, nn4397, nn4396, nn4395, nn4394, 
              nn4393, nn4392, nn4391} ), 
        .SUM( {\cal1_u132_XORCI_10|SUM_net , \cal1_u132_XORCI_9|SUM_net , 
              \cal1_u132_XORCI_8|SUM_net , \cal1_u132_XORCI_7|SUM_net , \cal1_u132_XORCI_6|SUM_net , 
              \cal1_u132_XORCI_5|SUM_net , \cal1_u132_XORCI_4|SUM_net , \cal1_u132_XORCI_3|SUM_net , 
              \cal1_u132_XORCI_2|SUM_net , \cal1_u132_XORCI_1|SUM_net , \cal1_u132_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4415 ( .DX(nn4415), .F0(dummy_36_), .F1(\cal1_u132_XORCI_10|SUM_net ), .F2(dummy_abc_3168_), .F3(dummy_abc_3169_) );
      defparam ii4415.CONFIG_DATA = 16'h8888;
      defparam ii4415.PLACE_LOCATION = "NONE";
      defparam ii4415.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4416 ( .DX(nn4416), .F0(dummy_36_), .F1(\cal1_u132_XORCI_1|SUM_net ), .F2(dummy_abc_3170_), .F3(dummy_abc_3171_) );
      defparam ii4416.CONFIG_DATA = 16'h8888;
      defparam ii4416.PLACE_LOCATION = "NONE";
      defparam ii4416.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4417 ( .DX(nn4417), .F0(dummy_36_), .F1(\cal1_u132_XORCI_2|SUM_net ), .F2(dummy_abc_3172_), .F3(dummy_abc_3173_) );
      defparam ii4417.CONFIG_DATA = 16'h8888;
      defparam ii4417.PLACE_LOCATION = "NONE";
      defparam ii4417.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4418 ( .DX(nn4418), .F0(dummy_36_), .F1(\cal1_u132_XORCI_3|SUM_net ), .F2(dummy_abc_3174_), .F3(dummy_abc_3175_) );
      defparam ii4418.CONFIG_DATA = 16'h8888;
      defparam ii4418.PLACE_LOCATION = "NONE";
      defparam ii4418.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4419 ( .DX(nn4419), .F0(dummy_36_), .F1(\cal1_u132_XORCI_4|SUM_net ), .F2(dummy_abc_3176_), .F3(dummy_abc_3177_) );
      defparam ii4419.CONFIG_DATA = 16'h8888;
      defparam ii4419.PLACE_LOCATION = "NONE";
      defparam ii4419.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4420 ( .DX(nn4420), .F0(dummy_36_), .F1(\cal1_u132_XORCI_5|SUM_net ), .F2(dummy_abc_3178_), .F3(dummy_abc_3179_) );
      defparam ii4420.CONFIG_DATA = 16'h8888;
      defparam ii4420.PLACE_LOCATION = "NONE";
      defparam ii4420.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4421 ( .DX(nn4421), .F0(dummy_36_), .F1(\cal1_u132_XORCI_6|SUM_net ), .F2(dummy_abc_3180_), .F3(dummy_abc_3181_) );
      defparam ii4421.CONFIG_DATA = 16'h8888;
      defparam ii4421.PLACE_LOCATION = "NONE";
      defparam ii4421.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4422 ( .DX(nn4422), .F0(dummy_36_), .F1(\cal1_u132_XORCI_7|SUM_net ), .F2(dummy_abc_3182_), .F3(dummy_abc_3183_) );
      defparam ii4422.CONFIG_DATA = 16'h8888;
      defparam ii4422.PLACE_LOCATION = "NONE";
      defparam ii4422.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4423 ( .DX(nn4423), .F0(dummy_36_), .F1(\cal1_u132_XORCI_8|SUM_net ), .F2(dummy_abc_3184_), .F3(dummy_abc_3185_) );
      defparam ii4423.CONFIG_DATA = 16'h8888;
      defparam ii4423.PLACE_LOCATION = "NONE";
      defparam ii4423.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4424 ( .DX(nn4424), .F0(dummy_36_), .F1(\cal1_u132_XORCI_9|SUM_net ), .F2(dummy_abc_3186_), .F3(dummy_abc_3187_) );
      defparam ii4424.CONFIG_DATA = 16'h8888;
      defparam ii4424.PLACE_LOCATION = "NONE";
      defparam ii4424.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4425 ( .DX(nn4425), .F0(en), .F1(iVsyn), .F2(\coefcal1_inEn__reg|Q_net ), .F3(\coefcal1_work__reg|Q_net ) );
      defparam ii4425.CONFIG_DATA = 16'hF8F0;
      defparam ii4425.PLACE_LOCATION = "NONE";
      defparam ii4425.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4426 ( .DX(nn4426), .F0(\a_mac_out[0]_coefcal1_u64_mac_0_ ), .F1(\a_mac_out[18]_coefcal1_u64_mac ), .F2(dummy_abc_3188_), .F3(dummy_abc_3189_) );
      defparam ii4426.CONFIG_DATA = 16'h6666;
      defparam ii4426.PLACE_LOCATION = "NONE";
      defparam ii4426.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4427 ( .DX(nn4427), .F0(\a_mac_out[0]_coefcal1_u64_mac_0_ ), .F1(\a_mac_out[18]_coefcal1_u64_mac ), .F2(dummy_abc_3190_), .F3(dummy_abc_3191_) );
      defparam ii4427.CONFIG_DATA = 16'h6666;
      defparam ii4427.PLACE_LOCATION = "NONE";
      defparam ii4427.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4428 ( .DX(nn4428), .F0(\a_mac_out[19]_coefcal1_u64_mac ), .F1(\a_mac_out[1]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_3192_), .F3(dummy_abc_3193_) );
      defparam ii4428.CONFIG_DATA = 16'h6666;
      defparam ii4428.PLACE_LOCATION = "NONE";
      defparam ii4428.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4429 ( .DX(nn4429), .F0(\a_mac_out[20]_coefcal1_u64_mac ), .F1(\a_mac_out[2]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_3194_), .F3(dummy_abc_3195_) );
      defparam ii4429.CONFIG_DATA = 16'h6666;
      defparam ii4429.PLACE_LOCATION = "NONE";
      defparam ii4429.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4430 ( .DX(nn4430), .F0(\a_mac_out[21]_coefcal1_u64_mac ), .F1(\a_mac_out[3]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_3196_), .F3(dummy_abc_3197_) );
      defparam ii4430.CONFIG_DATA = 16'h6666;
      defparam ii4430.PLACE_LOCATION = "NONE";
      defparam ii4430.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4431 ( .DX(nn4431), .F0(\a_mac_out[22]_coefcal1_u64_mac ), .F1(\a_mac_out[4]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_3198_), .F3(dummy_abc_3199_) );
      defparam ii4431.CONFIG_DATA = 16'h6666;
      defparam ii4431.PLACE_LOCATION = "NONE";
      defparam ii4431.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4432 ( .DX(nn4432), .F0(\a_mac_out[23]_coefcal1_u64_mac ), .F1(\a_mac_out[5]_coefcal1_u64_mac_0_ ), .F2(dummy_abc_3200_), .F3(dummy_abc_3201_) );
      defparam ii4432.CONFIG_DATA = 16'h6666;
      defparam ii4432.PLACE_LOCATION = "NONE";
      defparam ii4432.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4433 ( .DX(nn4433), .F0(\a_mac_out[6]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[0]_coefcal1_u64_mac ), .F2(dummy_abc_3202_), .F3(dummy_abc_3203_) );
      defparam ii4433.CONFIG_DATA = 16'h6666;
      defparam ii4433.PLACE_LOCATION = "NONE";
      defparam ii4433.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4434 ( .DX(nn4434), .F0(\a_mac_out[7]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[1]_coefcal1_u64_mac ), .F2(dummy_abc_3204_), .F3(dummy_abc_3205_) );
      defparam ii4434.CONFIG_DATA = 16'h6666;
      defparam ii4434.PLACE_LOCATION = "NONE";
      defparam ii4434.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4435 ( .DX(nn4435), .F0(\a_mac_out[8]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[2]_coefcal1_u64_mac ), .F2(dummy_abc_3206_), .F3(dummy_abc_3207_) );
      defparam ii4435.CONFIG_DATA = 16'h6666;
      defparam ii4435.PLACE_LOCATION = "NONE";
      defparam ii4435.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4436 ( .DX(nn4436), .F0(\a_mac_out[9]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[3]_coefcal1_u64_mac ), .F2(dummy_abc_3208_), .F3(dummy_abc_3209_) );
      defparam ii4436.CONFIG_DATA = 16'h6666;
      defparam ii4436.PLACE_LOCATION = "NONE";
      defparam ii4436.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4437 ( .DX(nn4437), .F0(\a_mac_out[10]_coefcal1_u64_mac_0_ ), .F1(\b_mac_out[4]_coefcal1_u64_mac ), .F2(dummy_abc_3210_), .F3(dummy_abc_3211_) );
      defparam ii4437.CONFIG_DATA = 16'h6666;
      defparam ii4437.PLACE_LOCATION = "NONE";
      defparam ii4437.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4438 ( .DX(nn4438), .F0(\a_mac_out[11]_coefcal1_u64_mac_0_ ), .F1(dummy_abc_3212_), .F2(dummy_abc_3213_), .F3(dummy_abc_3214_) );
      defparam ii4438.CONFIG_DATA = 16'hAAAA;
      defparam ii4438.PLACE_LOCATION = "NONE";
      defparam ii4438.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4439 ( .DX(nn4439), .F0(\a_mac_out[12]_coefcal1_u64_mac_0_ ), .F1(dummy_abc_3215_), .F2(dummy_abc_3216_), .F3(dummy_abc_3217_) );
      defparam ii4439.CONFIG_DATA = 16'hAAAA;
      defparam ii4439.PLACE_LOCATION = "NONE";
      defparam ii4439.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4440 ( .DX(nn4440), .F0(dummy_abc_3218_), .F1(dummy_abc_3219_), .F2(dummy_abc_3220_), .F3(dummy_abc_3221_) );
      defparam ii4440.CONFIG_DATA = 16'h0000;
      defparam ii4440.PLACE_LOCATION = "NONE";
      defparam ii4440.PCK_LOCATION = "NONE";
    scaler_ipc_adder_14 carry_14 ( 
        .CA( {a_acc_en_cal1_u137_mac, \a_mac_out[12]_coefcal1_u64_mac_0_ , 
              \a_mac_out[11]_coefcal1_u64_mac_0_ , \a_mac_out[10]_coefcal1_u64_mac_0_ , 
              \a_mac_out[9]_coefcal1_u64_mac_0_ , \a_mac_out[8]_coefcal1_u64_mac_0_ , 
              \a_mac_out[7]_coefcal1_u64_mac_0_ , \a_mac_out[6]_coefcal1_u64_mac_0_ , 
              \a_mac_out[5]_coefcal1_u64_mac_0_ , \a_mac_out[4]_coefcal1_u64_mac_0_ , 
              \a_mac_out[3]_coefcal1_u64_mac_0_ , \a_mac_out[2]_coefcal1_u64_mac_0_ , 
              \a_mac_out[1]_coefcal1_u64_mac_0_ , \a_mac_out[0]_coefcal1_u64_mac_0_ } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_137_ ), 
        .DX( {nn4440, nn4439, nn4438, nn4437, nn4436, nn4435, nn4434, nn4433, 
              nn4432, nn4431, nn4430, nn4429, nn4428, nn4427} ), 
        .SUM( {dummy_138_, \coefcal1_u64_XORCI_12|SUM_net , 
              \coefcal1_u64_XORCI_11|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , 
              \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u64_XORCI_8|SUM_net , 
              \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_6|SUM_net , 
              \coefcal1_u64_XORCI_5|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , 
              \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_2|SUM_net , 
              \coefcal1_u64_XORCI_1|SUM_net , \coefcal1_u64_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4457 ( .DX(nn4457), .F0(\a_mac_out[0]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[0]|Q_net ), .F2(dummy_abc_3222_), .F3(dummy_abc_3223_) );
      defparam ii4457.CONFIG_DATA = 16'h9999;
      defparam ii4457.PLACE_LOCATION = "NONE";
      defparam ii4457.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4458 ( .DX(nn4458), .F0(\a_mac_out[1]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[1]|Q_net ), .F2(dummy_abc_3224_), .F3(dummy_abc_3225_) );
      defparam ii4458.CONFIG_DATA = 16'h9999;
      defparam ii4458.PLACE_LOCATION = "NONE";
      defparam ii4458.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4459 ( .DX(nn4459), .F0(\a_mac_out[2]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[2]|Q_net ), .F2(dummy_abc_3226_), .F3(dummy_abc_3227_) );
      defparam ii4459.CONFIG_DATA = 16'h9999;
      defparam ii4459.PLACE_LOCATION = "NONE";
      defparam ii4459.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4460 ( .DX(nn4460), .F0(\a_mac_out[3]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[3]|Q_net ), .F2(dummy_abc_3228_), .F3(dummy_abc_3229_) );
      defparam ii4460.CONFIG_DATA = 16'h9999;
      defparam ii4460.PLACE_LOCATION = "NONE";
      defparam ii4460.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4461 ( .DX(nn4461), .F0(\a_mac_out[4]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[4]|Q_net ), .F2(dummy_abc_3230_), .F3(dummy_abc_3231_) );
      defparam ii4461.CONFIG_DATA = 16'h9999;
      defparam ii4461.PLACE_LOCATION = "NONE";
      defparam ii4461.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4462 ( .DX(nn4462), .F0(\a_mac_out[5]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[5]|Q_net ), .F2(dummy_abc_3232_), .F3(dummy_abc_3233_) );
      defparam ii4462.CONFIG_DATA = 16'h9999;
      defparam ii4462.PLACE_LOCATION = "NONE";
      defparam ii4462.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4463 ( .DX(nn4463), .F0(\a_mac_out[6]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[6]|Q_net ), .F2(dummy_abc_3234_), .F3(dummy_abc_3235_) );
      defparam ii4463.CONFIG_DATA = 16'h9999;
      defparam ii4463.PLACE_LOCATION = "NONE";
      defparam ii4463.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4464 ( .DX(nn4464), .F0(\a_mac_out[7]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[7]|Q_net ), .F2(dummy_abc_3236_), .F3(dummy_abc_3237_) );
      defparam ii4464.CONFIG_DATA = 16'h9999;
      defparam ii4464.PLACE_LOCATION = "NONE";
      defparam ii4464.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4465 ( .DX(nn4465), .F0(\a_mac_out[8]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[8]|Q_net ), .F2(dummy_abc_3238_), .F3(dummy_abc_3239_) );
      defparam ii4465.CONFIG_DATA = 16'h9999;
      defparam ii4465.PLACE_LOCATION = "NONE";
      defparam ii4465.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4466 ( .DX(nn4466), .F0(\a_mac_out[9]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[9]|Q_net ), .F2(dummy_abc_3240_), .F3(dummy_abc_3241_) );
      defparam ii4466.CONFIG_DATA = 16'h9999;
      defparam ii4466.PLACE_LOCATION = "NONE";
      defparam ii4466.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4467 ( .DX(nn4467), .F0(\a_mac_out[10]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[10]|Q_net ), .F2(dummy_abc_3242_), .F3(dummy_abc_3243_) );
      defparam ii4467.CONFIG_DATA = 16'h9999;
      defparam ii4467.PLACE_LOCATION = "NONE";
      defparam ii4467.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4468 ( .DX(nn4468), .F0(\a_mac_out[11]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[11]|Q_net ), .F2(dummy_abc_3244_), .F3(dummy_abc_3245_) );
      defparam ii4468.CONFIG_DATA = 16'h9999;
      defparam ii4468.PLACE_LOCATION = "NONE";
      defparam ii4468.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4469 ( .DX(nn4469), .F0(\a_mac_out[12]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[12]|Q_net ), .F2(dummy_abc_3246_), .F3(dummy_abc_3247_) );
      defparam ii4469.CONFIG_DATA = 16'h9999;
      defparam ii4469.PLACE_LOCATION = "NONE";
      defparam ii4469.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4470 ( .DX(nn4470), .F0(\a_mac_out[13]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[13]|Q_net ), .F2(dummy_abc_3248_), .F3(dummy_abc_3249_) );
      defparam ii4470.CONFIG_DATA = 16'h9999;
      defparam ii4470.PLACE_LOCATION = "NONE";
      defparam ii4470.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4471 ( .DX(nn4471), .F0(\a_mac_out[14]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[14]|Q_net ), .F2(dummy_abc_3250_), .F3(dummy_abc_3251_) );
      defparam ii4471.CONFIG_DATA = 16'h9999;
      defparam ii4471.PLACE_LOCATION = "NONE";
      defparam ii4471.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4472 ( .DX(nn4472), .F0(\a_mac_out[15]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[15]|Q_net ), .F2(dummy_abc_3252_), .F3(dummy_abc_3253_) );
      defparam ii4472.CONFIG_DATA = 16'h9999;
      defparam ii4472.PLACE_LOCATION = "NONE";
      defparam ii4472.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4473 ( .DX(nn4473), .F0(\a_mac_out[16]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[16]|Q_net ), .F2(dummy_abc_3254_), .F3(dummy_abc_3255_) );
      defparam ii4473.CONFIG_DATA = 16'h9999;
      defparam ii4473.PLACE_LOCATION = "NONE";
      defparam ii4473.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4474 ( .DX(nn4474), .F0(\a_mac_out[17]_coefcal1_u64_mac ), .F1(\coefcal1_working__reg[17]|Q_net ), .F2(dummy_abc_3256_), .F3(dummy_abc_3257_) );
      defparam ii4474.CONFIG_DATA = 16'h9999;
      defparam ii4474.PLACE_LOCATION = "NONE";
      defparam ii4474.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4475 ( .DX(nn4475), .F0(\coefcal1_working__reg[18]|Q_net ), .F1(nn4426), .F2(dummy_abc_3258_), .F3(dummy_abc_3259_) );
      defparam ii4475.CONFIG_DATA = 16'h9999;
      defparam ii4475.PLACE_LOCATION = "NONE";
      defparam ii4475.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4476 ( .DX(nn4476), .F0(\coefcal1_working__reg[19]|Q_net ), .F1(\coefcal1_u64_XORCI_1|SUM_net ), .F2(dummy_abc_3260_), .F3(dummy_abc_3261_) );
      defparam ii4476.CONFIG_DATA = 16'h9999;
      defparam ii4476.PLACE_LOCATION = "NONE";
      defparam ii4476.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4477 ( .DX(nn4477), .F0(\coefcal1_working__reg[20]|Q_net ), .F1(\coefcal1_u64_XORCI_2|SUM_net ), .F2(dummy_abc_3262_), .F3(dummy_abc_3263_) );
      defparam ii4477.CONFIG_DATA = 16'h9999;
      defparam ii4477.PLACE_LOCATION = "NONE";
      defparam ii4477.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4478 ( .DX(nn4478), .F0(\coefcal1_working__reg[21]|Q_net ), .F1(\coefcal1_u64_XORCI_3|SUM_net ), .F2(dummy_abc_3264_), .F3(dummy_abc_3265_) );
      defparam ii4478.CONFIG_DATA = 16'h9999;
      defparam ii4478.PLACE_LOCATION = "NONE";
      defparam ii4478.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4479 ( .DX(nn4479), .F0(\coefcal1_working__reg[22]|Q_net ), .F1(\coefcal1_u64_XORCI_4|SUM_net ), .F2(dummy_abc_3266_), .F3(dummy_abc_3267_) );
      defparam ii4479.CONFIG_DATA = 16'h9999;
      defparam ii4479.PLACE_LOCATION = "NONE";
      defparam ii4479.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4480 ( .DX(nn4480), .F0(\coefcal1_working__reg[23]|Q_net ), .F1(\coefcal1_u64_XORCI_5|SUM_net ), .F2(dummy_abc_3268_), .F3(dummy_abc_3269_) );
      defparam ii4480.CONFIG_DATA = 16'h9999;
      defparam ii4480.PLACE_LOCATION = "NONE";
      defparam ii4480.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4481 ( .DX(nn4481), .F0(\coefcal1_working__reg[24]|Q_net ), .F1(\coefcal1_u64_XORCI_6|SUM_net ), .F2(dummy_abc_3270_), .F3(dummy_abc_3271_) );
      defparam ii4481.CONFIG_DATA = 16'h9999;
      defparam ii4481.PLACE_LOCATION = "NONE";
      defparam ii4481.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4482 ( .DX(nn4482), .F0(\coefcal1_working__reg[25]|Q_net ), .F1(\coefcal1_u64_XORCI_7|SUM_net ), .F2(dummy_abc_3272_), .F3(dummy_abc_3273_) );
      defparam ii4482.CONFIG_DATA = 16'h9999;
      defparam ii4482.PLACE_LOCATION = "NONE";
      defparam ii4482.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4483 ( .DX(nn4483), .F0(\coefcal1_working__reg[26]|Q_net ), .F1(\coefcal1_u64_XORCI_8|SUM_net ), .F2(dummy_abc_3274_), .F3(dummy_abc_3275_) );
      defparam ii4483.CONFIG_DATA = 16'h9999;
      defparam ii4483.PLACE_LOCATION = "NONE";
      defparam ii4483.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4484 ( .DX(nn4484), .F0(\coefcal1_working__reg[27]|Q_net ), .F1(\coefcal1_u64_XORCI_9|SUM_net ), .F2(dummy_abc_3276_), .F3(dummy_abc_3277_) );
      defparam ii4484.CONFIG_DATA = 16'h9999;
      defparam ii4484.PLACE_LOCATION = "NONE";
      defparam ii4484.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4485 ( .DX(nn4485), .F0(\coefcal1_working__reg[28]|Q_net ), .F1(\coefcal1_u64_XORCI_10|SUM_net ), .F2(dummy_abc_3278_), .F3(dummy_abc_3279_) );
      defparam ii4485.CONFIG_DATA = 16'h9999;
      defparam ii4485.PLACE_LOCATION = "NONE";
      defparam ii4485.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4486 ( .DX(nn4486), .F0(\coefcal1_working__reg[29]|Q_net ), .F1(\coefcal1_u64_XORCI_11|SUM_net ), .F2(dummy_abc_3280_), .F3(dummy_abc_3281_) );
      defparam ii4486.CONFIG_DATA = 16'h9999;
      defparam ii4486.PLACE_LOCATION = "NONE";
      defparam ii4486.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4487 ( .DX(nn4487), .F0(\coefcal1_working__reg[30]|Q_net ), .F1(\coefcal1_u64_XORCI_12|SUM_net ), .F2(dummy_abc_3282_), .F3(dummy_abc_3283_) );
      defparam ii4487.CONFIG_DATA = 16'h9999;
      defparam ii4487.PLACE_LOCATION = "NONE";
      defparam ii4487.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4488 ( .DX(nn4488), .F0(\coefcal1_working__reg[31]|Q_net ), .F1(dummy_abc_3284_), .F2(dummy_abc_3285_), .F3(dummy_abc_3286_) );
      defparam ii4488.CONFIG_DATA = 16'h5555;
      defparam ii4488.PLACE_LOCATION = "NONE";
      defparam ii4488.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4489 ( .DX(nn4489), .F0(\coefcal1_working__reg[32]|Q_net ), .F1(dummy_abc_3287_), .F2(dummy_abc_3288_), .F3(dummy_abc_3289_) );
      defparam ii4489.CONFIG_DATA = 16'h5555;
      defparam ii4489.PLACE_LOCATION = "NONE";
      defparam ii4489.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4490 ( .DX(nn4490), .F0(dummy_abc_3290_), .F1(dummy_abc_3291_), .F2(dummy_abc_3292_), .F3(dummy_abc_3293_) );
      defparam ii4490.CONFIG_DATA = 16'hFFFF;
      defparam ii4490.PLACE_LOCATION = "NONE";
      defparam ii4490.PCK_LOCATION = "NONE";
    scaler_ipc_adder_34 carry_34 ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, \coefcal1_u64_XORCI_12|SUM_net , 
              \coefcal1_u64_XORCI_11|SUM_net , \coefcal1_u64_XORCI_10|SUM_net , 
              \coefcal1_u64_XORCI_9|SUM_net , \coefcal1_u64_XORCI_8|SUM_net , 
              \coefcal1_u64_XORCI_7|SUM_net , \coefcal1_u64_XORCI_6|SUM_net , 
              \coefcal1_u64_XORCI_5|SUM_net , \coefcal1_u64_XORCI_4|SUM_net , 
              \coefcal1_u64_XORCI_3|SUM_net , \coefcal1_u64_XORCI_2|SUM_net , 
              \coefcal1_u64_XORCI_1|SUM_net , nn4426, \a_mac_out[17]_coefcal1_u64_mac , 
              \a_mac_out[16]_coefcal1_u64_mac , \a_mac_out[15]_coefcal1_u64_mac , 
              \a_mac_out[14]_coefcal1_u64_mac , \a_mac_out[13]_coefcal1_u64_mac , 
              \a_mac_out[12]_coefcal1_u64_mac , \a_mac_out[11]_coefcal1_u64_mac , 
              \a_mac_out[10]_coefcal1_u64_mac , \a_mac_out[9]_coefcal1_u64_mac , 
              \a_mac_out[8]_coefcal1_u64_mac , \a_mac_out[7]_coefcal1_u64_mac , 
              \a_mac_out[6]_coefcal1_u64_mac , \a_mac_out[5]_coefcal1_u64_mac , 
              \a_mac_out[4]_coefcal1_u64_mac , \a_mac_out[3]_coefcal1_u64_mac , 
              \a_mac_out[2]_coefcal1_u64_mac , \a_mac_out[1]_coefcal1_u64_mac , 
              \a_mac_out[0]_coefcal1_u64_mac } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_850_ ), 
        .DX( {nn4490, nn4489, nn4488, nn4487, nn4486, nn4485, nn4484, nn4483, 
              nn4482, nn4481, nn4480, nn4479, nn4478, nn4477, nn4476, nn4475, 
              nn4474, nn4473, nn4472, nn4471, nn4470, nn4469, nn4468, nn4467, 
              nn4466, nn4465, nn4464, nn4463, nn4462, nn4461, nn4460, nn4459, 
              nn4458, nn4457} ), 
        .SUM( {\coefcal1_u8_XORCI_33|SUM_net , dummy_851_, dummy_852_, dummy_853_, 
              dummy_854_, dummy_855_, dummy_856_, dummy_857_, dummy_858_, dummy_859_, 
              dummy_860_, dummy_861_, dummy_862_, dummy_863_, dummy_864_, dummy_865_, 
              dummy_866_, dummy_867_, dummy_868_, dummy_869_, dummy_870_, dummy_871_, 
              dummy_872_, dummy_873_, dummy_874_, dummy_875_, dummy_876_, dummy_877_, 
              dummy_878_, dummy_879_, dummy_880_, dummy_881_, dummy_882_, dummy_883_} )
      );
    CS_LUT4_PRIM ii4527 ( .DX(nn4527), .F0(dummy_850_), .F1(dummy_abc_3294_), .F2(dummy_abc_3295_), .F3(dummy_abc_3296_) );
      defparam ii4527.CONFIG_DATA = 16'h5555;
      defparam ii4527.PLACE_LOCATION = "NONE";
      defparam ii4527.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4528 ( .DX(nn4528), .F0(nn0886), .F1(dummy_abc_3297_), .F2(dummy_abc_3298_), .F3(dummy_abc_3299_) );
      defparam ii4528.CONFIG_DATA = 16'h5555;
      defparam ii4528.PLACE_LOCATION = "NONE";
      defparam ii4528.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4529 ( .DX(nn4529), .F0(\u2_XORCI_1|SUM_net ), .F1(dummy_abc_3300_), .F2(dummy_abc_3301_), .F3(dummy_abc_3302_) );
      defparam ii4529.CONFIG_DATA = 16'hAAAA;
      defparam ii4529.PLACE_LOCATION = "NONE";
      defparam ii4529.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4530 ( .DX(nn4530), .F0(\u2_XORCI_2|SUM_net ), .F1(dummy_abc_3303_), .F2(dummy_abc_3304_), .F3(dummy_abc_3305_) );
      defparam ii4530.CONFIG_DATA = 16'hAAAA;
      defparam ii4530.PLACE_LOCATION = "NONE";
      defparam ii4530.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4531 ( .DX(nn4531), .F0(\u2_XORCI_3|SUM_net ), .F1(dummy_abc_3306_), .F2(dummy_abc_3307_), .F3(dummy_abc_3308_) );
      defparam ii4531.CONFIG_DATA = 16'hAAAA;
      defparam ii4531.PLACE_LOCATION = "NONE";
      defparam ii4531.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4532 ( .DX(nn4532), .F0(\u2_XORCI_4|SUM_net ), .F1(dummy_abc_3309_), .F2(dummy_abc_3310_), .F3(dummy_abc_3311_) );
      defparam ii4532.CONFIG_DATA = 16'hAAAA;
      defparam ii4532.PLACE_LOCATION = "NONE";
      defparam ii4532.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4533 ( .DX(nn4533), .F0(\u2_XORCI_5|SUM_net ), .F1(dummy_abc_3312_), .F2(dummy_abc_3313_), .F3(dummy_abc_3314_) );
      defparam ii4533.CONFIG_DATA = 16'hAAAA;
      defparam ii4533.PLACE_LOCATION = "NONE";
      defparam ii4533.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4534 ( .DX(nn4534), .F0(\u2_XORCI_6|SUM_net ), .F1(dummy_abc_3315_), .F2(dummy_abc_3316_), .F3(dummy_abc_3317_) );
      defparam ii4534.CONFIG_DATA = 16'hAAAA;
      defparam ii4534.PLACE_LOCATION = "NONE";
      defparam ii4534.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4535 ( .DX(nn4535), .F0(\u2_XORCI_7|SUM_net ), .F1(dummy_abc_3318_), .F2(dummy_abc_3319_), .F3(dummy_abc_3320_) );
      defparam ii4535.CONFIG_DATA = 16'hAAAA;
      defparam ii4535.PLACE_LOCATION = "NONE";
      defparam ii4535.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4536 ( .DX(nn4536), .F0(\u2_XORCI_8|SUM_net ), .F1(dummy_abc_3321_), .F2(dummy_abc_3322_), .F3(dummy_abc_3323_) );
      defparam ii4536.CONFIG_DATA = 16'hAAAA;
      defparam ii4536.PLACE_LOCATION = "NONE";
      defparam ii4536.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4537 ( .DX(nn4537), .F0(\u2_XORCI_9|SUM_net ), .F1(dummy_abc_3324_), .F2(dummy_abc_3325_), .F3(dummy_abc_3326_) );
      defparam ii4537.CONFIG_DATA = 16'hAAAA;
      defparam ii4537.PLACE_LOCATION = "NONE";
      defparam ii4537.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4538 ( .DX(nn4538), .F0(\u2_XORCI_10|SUM_net ), .F1(dummy_abc_3327_), .F2(dummy_abc_3328_), .F3(dummy_abc_3329_) );
      defparam ii4538.CONFIG_DATA = 16'hAAAA;
      defparam ii4538.PLACE_LOCATION = "NONE";
      defparam ii4538.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_277_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_dinxy_cen_cal1_u137_mac} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_17_ ), 
        .DX( {nn4538, nn4537, nn4536, nn4535, nn4534, nn4533, nn4532, nn4531, 
              nn4530, nn4529, nn4528} ), 
        .SUM( {\coefcal1_u59_XORCI_10|SUM_net , \coefcal1_u59_XORCI_9|SUM_net , 
              \coefcal1_u59_XORCI_8|SUM_net , \coefcal1_u59_XORCI_7|SUM_net , 
              \coefcal1_u59_XORCI_6|SUM_net , \coefcal1_u59_XORCI_5|SUM_net , 
              \coefcal1_u59_XORCI_4|SUM_net , \coefcal1_u59_XORCI_3|SUM_net , 
              \coefcal1_u59_XORCI_2|SUM_net , \coefcal1_u59_XORCI_1|SUM_net , 
              \coefcal1_u59_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4552 ( .DX(nn4552), .F0(nn0886), .F1(dummy_abc_3330_), .F2(dummy_abc_3331_), .F3(dummy_abc_3332_) );
      defparam ii4552.CONFIG_DATA = 16'h5555;
      defparam ii4552.PLACE_LOCATION = "NONE";
      defparam ii4552.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4553 ( .DX(nn4553), .F0(\u3_XORCI_1|SUM_net ), .F1(dummy_abc_3333_), .F2(dummy_abc_3334_), .F3(dummy_abc_3335_) );
      defparam ii4553.CONFIG_DATA = 16'h5555;
      defparam ii4553.PLACE_LOCATION = "NONE";
      defparam ii4553.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4554 ( .DX(nn4554), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3336_), .F3(dummy_abc_3337_) );
      defparam ii4554.CONFIG_DATA = 16'h9999;
      defparam ii4554.PLACE_LOCATION = "NONE";
      defparam ii4554.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4555 ( .DX(nn4555), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3338_), .F3(dummy_abc_3339_) );
      defparam ii4555.CONFIG_DATA = 16'h9999;
      defparam ii4555.PLACE_LOCATION = "NONE";
      defparam ii4555.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4556 ( .DX(nn4556), .F0(yBgn[1]), .F1(yEnd[1]), .F2(dummy_abc_3340_), .F3(dummy_abc_3341_) );
      defparam ii4556.CONFIG_DATA = 16'h9999;
      defparam ii4556.PLACE_LOCATION = "NONE";
      defparam ii4556.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4557 ( .DX(nn4557), .F0(yBgn[2]), .F1(yEnd[2]), .F2(dummy_abc_3342_), .F3(dummy_abc_3343_) );
      defparam ii4557.CONFIG_DATA = 16'h9999;
      defparam ii4557.PLACE_LOCATION = "NONE";
      defparam ii4557.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4558 ( .DX(nn4558), .F0(yBgn[3]), .F1(yEnd[3]), .F2(dummy_abc_3344_), .F3(dummy_abc_3345_) );
      defparam ii4558.CONFIG_DATA = 16'h9999;
      defparam ii4558.PLACE_LOCATION = "NONE";
      defparam ii4558.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4559 ( .DX(nn4559), .F0(yBgn[4]), .F1(yEnd[4]), .F2(dummy_abc_3346_), .F3(dummy_abc_3347_) );
      defparam ii4559.CONFIG_DATA = 16'h9999;
      defparam ii4559.PLACE_LOCATION = "NONE";
      defparam ii4559.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4560 ( .DX(nn4560), .F0(yBgn[5]), .F1(yEnd[5]), .F2(dummy_abc_3348_), .F3(dummy_abc_3349_) );
      defparam ii4560.CONFIG_DATA = 16'h9999;
      defparam ii4560.PLACE_LOCATION = "NONE";
      defparam ii4560.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4561 ( .DX(nn4561), .F0(yBgn[6]), .F1(yEnd[6]), .F2(dummy_abc_3350_), .F3(dummy_abc_3351_) );
      defparam ii4561.CONFIG_DATA = 16'h9999;
      defparam ii4561.PLACE_LOCATION = "NONE";
      defparam ii4561.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4562 ( .DX(nn4562), .F0(yBgn[7]), .F1(yEnd[7]), .F2(dummy_abc_3352_), .F3(dummy_abc_3353_) );
      defparam ii4562.CONFIG_DATA = 16'h9999;
      defparam ii4562.PLACE_LOCATION = "NONE";
      defparam ii4562.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4563 ( .DX(nn4563), .F0(yBgn[8]), .F1(yEnd[8]), .F2(dummy_abc_3354_), .F3(dummy_abc_3355_) );
      defparam ii4563.CONFIG_DATA = 16'h9999;
      defparam ii4563.PLACE_LOCATION = "NONE";
      defparam ii4563.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4564 ( .DX(nn4564), .F0(yBgn[9]), .F1(yEnd[9]), .F2(dummy_abc_3356_), .F3(dummy_abc_3357_) );
      defparam ii4564.CONFIG_DATA = 16'h9999;
      defparam ii4564.PLACE_LOCATION = "NONE";
      defparam ii4564.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4565 ( .DX(nn4565), .F0(yBgn[10]), .F1(yEnd[10]), .F2(dummy_abc_3358_), .F3(dummy_abc_3359_) );
      defparam ii4565.CONFIG_DATA = 16'h9999;
      defparam ii4565.PLACE_LOCATION = "NONE";
      defparam ii4565.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4566 ( .DX(nn4566), .F0(dummy_abc_3360_), .F1(dummy_abc_3361_), .F2(dummy_abc_3362_), .F3(dummy_abc_3363_) );
      defparam ii4566.CONFIG_DATA = 16'hFFFF;
      defparam ii4566.PLACE_LOCATION = "NONE";
      defparam ii4566.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_281_ ( 
        .CA( {a_acc_en_cal1_u137_mac, yEnd[10], yEnd[9], yEnd[8], yEnd[7], 
              yEnd[6], yEnd[5], yEnd[4], yEnd[3], yEnd[2], yEnd[1], yEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_76_ ), 
        .DX( {nn4566, nn4565, nn4564, nn4563, nn4562, nn4561, nn4560, nn4559, 
              nn4558, nn4557, nn4556, nn4555} ), 
        .SUM( {dummy_77_, \coefcal1_u7_XORCI_10|SUM_net , 
              \coefcal1_u7_XORCI_9|SUM_net , \coefcal1_u7_XORCI_8|SUM_net , 
              \coefcal1_u7_XORCI_7|SUM_net , \coefcal1_u7_XORCI_6|SUM_net , 
              \coefcal1_u7_XORCI_5|SUM_net , \coefcal1_u7_XORCI_4|SUM_net , 
              \coefcal1_u7_XORCI_3|SUM_net , \coefcal1_u7_XORCI_2|SUM_net , 
              \coefcal1_u7_XORCI_1|SUM_net , \coefcal1_u7_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4581 ( .DX(nn4581), .F0(\coefcal1_u7_XORCI_1|SUM_net ), .F1(dummy_abc_3364_), .F2(dummy_abc_3365_), .F3(dummy_abc_3366_) );
      defparam ii4581.CONFIG_DATA = 16'hAAAA;
      defparam ii4581.PLACE_LOCATION = "NONE";
      defparam ii4581.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4582 ( .DX(nn4582), .F0(\coefcal1_u7_XORCI_2|SUM_net ), .F1(dummy_abc_3367_), .F2(dummy_abc_3368_), .F3(dummy_abc_3369_) );
      defparam ii4582.CONFIG_DATA = 16'hAAAA;
      defparam ii4582.PLACE_LOCATION = "NONE";
      defparam ii4582.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4583 ( .DX(nn4583), .F0(\coefcal1_u7_XORCI_3|SUM_net ), .F1(dummy_abc_3370_), .F2(dummy_abc_3371_), .F3(dummy_abc_3372_) );
      defparam ii4583.CONFIG_DATA = 16'hAAAA;
      defparam ii4583.PLACE_LOCATION = "NONE";
      defparam ii4583.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4584 ( .DX(nn4584), .F0(\coefcal1_u7_XORCI_4|SUM_net ), .F1(dummy_abc_3373_), .F2(dummy_abc_3374_), .F3(dummy_abc_3375_) );
      defparam ii4584.CONFIG_DATA = 16'hAAAA;
      defparam ii4584.PLACE_LOCATION = "NONE";
      defparam ii4584.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4585 ( .DX(nn4585), .F0(\coefcal1_u7_XORCI_5|SUM_net ), .F1(dummy_abc_3376_), .F2(dummy_abc_3377_), .F3(dummy_abc_3378_) );
      defparam ii4585.CONFIG_DATA = 16'hAAAA;
      defparam ii4585.PLACE_LOCATION = "NONE";
      defparam ii4585.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4586 ( .DX(nn4586), .F0(\coefcal1_u7_XORCI_6|SUM_net ), .F1(dummy_abc_3379_), .F2(dummy_abc_3380_), .F3(dummy_abc_3381_) );
      defparam ii4586.CONFIG_DATA = 16'hAAAA;
      defparam ii4586.PLACE_LOCATION = "NONE";
      defparam ii4586.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4587 ( .DX(nn4587), .F0(\coefcal1_u7_XORCI_7|SUM_net ), .F1(dummy_abc_3382_), .F2(dummy_abc_3383_), .F3(dummy_abc_3384_) );
      defparam ii4587.CONFIG_DATA = 16'hAAAA;
      defparam ii4587.PLACE_LOCATION = "NONE";
      defparam ii4587.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4588 ( .DX(nn4588), .F0(\coefcal1_u7_XORCI_8|SUM_net ), .F1(dummy_abc_3385_), .F2(dummy_abc_3386_), .F3(dummy_abc_3387_) );
      defparam ii4588.CONFIG_DATA = 16'hAAAA;
      defparam ii4588.PLACE_LOCATION = "NONE";
      defparam ii4588.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4589 ( .DX(nn4589), .F0(\coefcal1_u7_XORCI_9|SUM_net ), .F1(dummy_abc_3388_), .F2(dummy_abc_3389_), .F3(dummy_abc_3390_) );
      defparam ii4589.CONFIG_DATA = 16'hAAAA;
      defparam ii4589.PLACE_LOCATION = "NONE";
      defparam ii4589.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4590 ( .DX(nn4590), .F0(\coefcal1_u7_XORCI_10|SUM_net ), .F1(dummy_abc_3391_), .F2(dummy_abc_3392_), .F3(dummy_abc_3393_) );
      defparam ii4590.CONFIG_DATA = 16'hAAAA;
      defparam ii4590.PLACE_LOCATION = "NONE";
      defparam ii4590.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_278_ ( 
        .CA( {a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, 
              a_acc_en_cal1_u137_mac, a_acc_en_cal1_u137_mac, a_dinxy_cen_cal1_u137_mac} ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_18_ ), 
        .DX( {nn4590, nn4589, nn4588, nn4587, nn4586, nn4585, nn4584, nn4583, 
              nn4582, nn4581, nn4554} ), 
        .SUM( {\coefcal1_u60_XORCI_10|SUM_net , \coefcal1_u60_XORCI_9|SUM_net , 
              \coefcal1_u60_XORCI_8|SUM_net , \coefcal1_u60_XORCI_7|SUM_net , 
              \coefcal1_u60_XORCI_6|SUM_net , \coefcal1_u60_XORCI_5|SUM_net , 
              \coefcal1_u60_XORCI_4|SUM_net , \coefcal1_u60_XORCI_3|SUM_net , 
              \coefcal1_u60_XORCI_2|SUM_net , \coefcal1_u60_XORCI_1|SUM_net , 
              \coefcal1_u60_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4604 ( .DX(nn4604), .F0(yBgn[0]), .F1(yEnd[0]), .F2(dummy_abc_3394_), .F3(dummy_abc_3395_) );
      defparam ii4604.CONFIG_DATA = 16'h9999;
      defparam ii4604.PLACE_LOCATION = "NONE";
      defparam ii4604.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4605 ( .DX(nn4605), .F0(dIn[0]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3396_) );
      defparam ii4605.CONFIG_DATA = 16'h0202;
      defparam ii4605.PLACE_LOCATION = "NONE";
      defparam ii4605.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4606 ( .DX(nn4606), .F0(\inputctrl1_xAddress__reg[1]|Q_net ), .F1(\inputctrl1_xAddress__reg[5]|Q_net ), .F2(\inputctrl1_xCal__reg[11]|Q_net ), .F3(\inputctrl1_xCal__reg[7]|Q_net ) );
      defparam ii4606.CONFIG_DATA = 16'h8241;
      defparam ii4606.PLACE_LOCATION = "NONE";
      defparam ii4606.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4607 ( .DX(nn4607), .F0(\inputctrl1_xAddress__reg[7]|Q_net ), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(\inputctrl1_xCal__reg[13]|Q_net ), .F3(\inputctrl1_xCal__reg[15]|Q_net ) );
      defparam ii4607.CONFIG_DATA = 16'h8421;
      defparam ii4607.PLACE_LOCATION = "NONE";
      defparam ii4607.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4608 ( .DX(nn4608), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(\inputctrl1_xAddress__reg[3]|Q_net ), .F2(\inputctrl1_xCal__reg[6]|Q_net ), .F3(\inputctrl1_xCal__reg[9]|Q_net ) );
      defparam ii4608.CONFIG_DATA = 16'h8421;
      defparam ii4608.PLACE_LOCATION = "NONE";
      defparam ii4608.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4609 ( .DX(nn4609), .F0(\inputctrl1_xAddress__reg[2]|Q_net ), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(\inputctrl1_xCal__reg[12]|Q_net ), .F3(\inputctrl1_xCal__reg[8]|Q_net ) );
      defparam ii4609.CONFIG_DATA = 16'h8241;
      defparam ii4609.PLACE_LOCATION = "NONE";
      defparam ii4609.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4610 ( .DX(nn4610), .F0(\inputctrl1_xAddress__reg[10]|Q_net ), .F1(\inputctrl1_xAddress__reg[4]|Q_net ), .F2(\inputctrl1_xCal__reg[10]|Q_net ), .F3(\inputctrl1_xCal__reg[16]|Q_net ) );
      defparam ii4610.CONFIG_DATA = 16'h8241;
      defparam ii4610.PLACE_LOCATION = "NONE";
      defparam ii4610.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4611 ( .DX(nn4611), .F0(nn4607), .F1(nn4608), .F2(nn4609), .F3(nn4610) );
      defparam ii4611.CONFIG_DATA = 16'h8000;
      defparam ii4611.PLACE_LOCATION = "NONE";
      defparam ii4611.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4612 ( .DX(nn4612), .F0(\inputctrl1_xAddress__reg[8]|Q_net ), .F1(\inputctrl1_xCal__reg[14]|Q_net ), .F2(nn4606), .F3(nn4611) );
      defparam ii4612.CONFIG_DATA = 16'h9000;
      defparam ii4612.PLACE_LOCATION = "NONE";
      defparam ii4612.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4613 ( .DX(nn4613), .F0(yBgn[0]), .F1(\inputctrl1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_3397_), .F3(dummy_abc_3398_) );
      defparam ii4613.CONFIG_DATA = 16'h9999;
      defparam ii4613.PLACE_LOCATION = "NONE";
      defparam ii4613.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4614 ( .DX(nn4614), .F0(yBgn[1]), .F1(\inputctrl1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_3399_), .F3(dummy_abc_3400_) );
      defparam ii4614.CONFIG_DATA = 16'h9999;
      defparam ii4614.PLACE_LOCATION = "NONE";
      defparam ii4614.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4615 ( .DX(nn4615), .F0(yBgn[2]), .F1(\inputctrl1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_3401_), .F3(dummy_abc_3402_) );
      defparam ii4615.CONFIG_DATA = 16'h9999;
      defparam ii4615.PLACE_LOCATION = "NONE";
      defparam ii4615.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4616 ( .DX(nn4616), .F0(yBgn[3]), .F1(\inputctrl1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_3403_), .F3(dummy_abc_3404_) );
      defparam ii4616.CONFIG_DATA = 16'h9999;
      defparam ii4616.PLACE_LOCATION = "NONE";
      defparam ii4616.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4617 ( .DX(nn4617), .F0(yBgn[4]), .F1(\inputctrl1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_3405_), .F3(dummy_abc_3406_) );
      defparam ii4617.CONFIG_DATA = 16'h9999;
      defparam ii4617.PLACE_LOCATION = "NONE";
      defparam ii4617.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4618 ( .DX(nn4618), .F0(yBgn[5]), .F1(\inputctrl1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_3407_), .F3(dummy_abc_3408_) );
      defparam ii4618.CONFIG_DATA = 16'h9999;
      defparam ii4618.PLACE_LOCATION = "NONE";
      defparam ii4618.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4619 ( .DX(nn4619), .F0(yBgn[6]), .F1(\inputctrl1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_3409_), .F3(dummy_abc_3410_) );
      defparam ii4619.CONFIG_DATA = 16'h9999;
      defparam ii4619.PLACE_LOCATION = "NONE";
      defparam ii4619.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4620 ( .DX(nn4620), .F0(yBgn[7]), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_3411_), .F3(dummy_abc_3412_) );
      defparam ii4620.CONFIG_DATA = 16'h9999;
      defparam ii4620.PLACE_LOCATION = "NONE";
      defparam ii4620.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4621 ( .DX(nn4621), .F0(yBgn[8]), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_3413_), .F3(dummy_abc_3414_) );
      defparam ii4621.CONFIG_DATA = 16'h9999;
      defparam ii4621.PLACE_LOCATION = "NONE";
      defparam ii4621.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4622 ( .DX(nn4622), .F0(yBgn[9]), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_3415_), .F3(dummy_abc_3416_) );
      defparam ii4622.CONFIG_DATA = 16'h9999;
      defparam ii4622.PLACE_LOCATION = "NONE";
      defparam ii4622.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4623 ( .DX(nn4623), .F0(yBgn[10]), .F1(\inputctrl1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_3417_), .F3(dummy_abc_3418_) );
      defparam ii4623.CONFIG_DATA = 16'h9999;
      defparam ii4623.PLACE_LOCATION = "NONE";
      defparam ii4623.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4624 ( .DX(nn4624), .F0(dummy_abc_3419_), .F1(dummy_abc_3420_), .F2(dummy_abc_3421_), .F3(dummy_abc_3422_) );
      defparam ii4624.CONFIG_DATA = 16'hFFFF;
      defparam ii4624.PLACE_LOCATION = "NONE";
      defparam ii4624.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_288_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \inputctrl1_yAddress__reg[10]|Q_net , 
              \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net , 
              \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net , 
              \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net , 
              \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net , 
              \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_92_ ), 
        .DX( {nn4624, nn4623, nn4622, nn4621, nn4620, nn4619, nn4618, nn4617, 
              nn4616, nn4615, nn4614, nn4613} ), 
        .SUM( {\inputctrl1_u39_XORCI_11|SUM_net , dummy_93_, dummy_94_, dummy_95_, 
              dummy_96_, dummy_97_, dummy_98_, dummy_99_, dummy_100_, dummy_101_, 
              dummy_102_, dummy_103_} )
      );
    CS_LUT4_PRIM ii4639 ( .DX(nn4639), .F0(\inputctrl1_yAddress__reg[2]|Q_net ), .F1(\inputctrl1_yAddress__reg[6]|Q_net ), .F2(\inputctrl1_yCal__reg[12]|Q_net ), .F3(\inputctrl1_yCal__reg[8]|Q_net ) );
      defparam ii4639.CONFIG_DATA = 16'h8241;
      defparam ii4639.PLACE_LOCATION = "NONE";
      defparam ii4639.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4640 ( .DX(nn4640), .F0(\inputctrl1_yAddress__reg[10]|Q_net ), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(\inputctrl1_yCal__reg[14]|Q_net ), .F3(\inputctrl1_yCal__reg[16]|Q_net ) );
      defparam ii4640.CONFIG_DATA = 16'h8241;
      defparam ii4640.PLACE_LOCATION = "NONE";
      defparam ii4640.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4641 ( .DX(nn4641), .F0(\inputctrl1_yAddress__reg[3]|Q_net ), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(\inputctrl1_yCal__reg[13]|Q_net ), .F3(\inputctrl1_yCal__reg[9]|Q_net ) );
      defparam ii4641.CONFIG_DATA = 16'h8241;
      defparam ii4641.PLACE_LOCATION = "NONE";
      defparam ii4641.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4642 ( .DX(nn4642), .F0(\inputctrl1_yAddress__reg[1]|Q_net ), .F1(\inputctrl1_yAddress__reg[5]|Q_net ), .F2(\inputctrl1_yCal__reg[11]|Q_net ), .F3(\inputctrl1_yCal__reg[7]|Q_net ) );
      defparam ii4642.CONFIG_DATA = 16'h8241;
      defparam ii4642.PLACE_LOCATION = "NONE";
      defparam ii4642.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4643 ( .DX(nn4643), .F0(\inputctrl1_yAddress__reg[4]|Q_net ), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(\inputctrl1_yCal__reg[10]|Q_net ), .F3(\inputctrl1_yCal__reg[15]|Q_net ) );
      defparam ii4643.CONFIG_DATA = 16'h8421;
      defparam ii4643.PLACE_LOCATION = "NONE";
      defparam ii4643.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4644 ( .DX(nn4644), .F0(nn4640), .F1(nn4641), .F2(nn4642), .F3(nn4643) );
      defparam ii4644.CONFIG_DATA = 16'h8000;
      defparam ii4644.PLACE_LOCATION = "NONE";
      defparam ii4644.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4645 ( .DX(nn4645), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(\inputctrl1_yCal__reg[6]|Q_net ), .F2(nn4639), .F3(nn4644) );
      defparam ii4645.CONFIG_DATA = 16'h9000;
      defparam ii4645.PLACE_LOCATION = "NONE";
      defparam ii4645.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4646 ( .DX(nn4646), .F0(yEnd[0]), .F1(\inputctrl1_yAddress__reg[0]|Q_net ), .F2(dummy_abc_3423_), .F3(dummy_abc_3424_) );
      defparam ii4646.CONFIG_DATA = 16'h9999;
      defparam ii4646.PLACE_LOCATION = "NONE";
      defparam ii4646.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4647 ( .DX(nn4647), .F0(yEnd[1]), .F1(\inputctrl1_yAddress__reg[1]|Q_net ), .F2(dummy_abc_3425_), .F3(dummy_abc_3426_) );
      defparam ii4647.CONFIG_DATA = 16'h9999;
      defparam ii4647.PLACE_LOCATION = "NONE";
      defparam ii4647.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4648 ( .DX(nn4648), .F0(yEnd[2]), .F1(\inputctrl1_yAddress__reg[2]|Q_net ), .F2(dummy_abc_3427_), .F3(dummy_abc_3428_) );
      defparam ii4648.CONFIG_DATA = 16'h9999;
      defparam ii4648.PLACE_LOCATION = "NONE";
      defparam ii4648.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4649 ( .DX(nn4649), .F0(yEnd[3]), .F1(\inputctrl1_yAddress__reg[3]|Q_net ), .F2(dummy_abc_3429_), .F3(dummy_abc_3430_) );
      defparam ii4649.CONFIG_DATA = 16'h9999;
      defparam ii4649.PLACE_LOCATION = "NONE";
      defparam ii4649.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4650 ( .DX(nn4650), .F0(yEnd[4]), .F1(\inputctrl1_yAddress__reg[4]|Q_net ), .F2(dummy_abc_3431_), .F3(dummy_abc_3432_) );
      defparam ii4650.CONFIG_DATA = 16'h9999;
      defparam ii4650.PLACE_LOCATION = "NONE";
      defparam ii4650.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4651 ( .DX(nn4651), .F0(yEnd[5]), .F1(\inputctrl1_yAddress__reg[5]|Q_net ), .F2(dummy_abc_3433_), .F3(dummy_abc_3434_) );
      defparam ii4651.CONFIG_DATA = 16'h9999;
      defparam ii4651.PLACE_LOCATION = "NONE";
      defparam ii4651.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4652 ( .DX(nn4652), .F0(yEnd[6]), .F1(\inputctrl1_yAddress__reg[6]|Q_net ), .F2(dummy_abc_3435_), .F3(dummy_abc_3436_) );
      defparam ii4652.CONFIG_DATA = 16'h9999;
      defparam ii4652.PLACE_LOCATION = "NONE";
      defparam ii4652.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4653 ( .DX(nn4653), .F0(yEnd[7]), .F1(\inputctrl1_yAddress__reg[7]|Q_net ), .F2(dummy_abc_3437_), .F3(dummy_abc_3438_) );
      defparam ii4653.CONFIG_DATA = 16'h9999;
      defparam ii4653.PLACE_LOCATION = "NONE";
      defparam ii4653.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4654 ( .DX(nn4654), .F0(yEnd[8]), .F1(\inputctrl1_yAddress__reg[8]|Q_net ), .F2(dummy_abc_3439_), .F3(dummy_abc_3440_) );
      defparam ii4654.CONFIG_DATA = 16'h9999;
      defparam ii4654.PLACE_LOCATION = "NONE";
      defparam ii4654.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4655 ( .DX(nn4655), .F0(yEnd[9]), .F1(\inputctrl1_yAddress__reg[9]|Q_net ), .F2(dummy_abc_3441_), .F3(dummy_abc_3442_) );
      defparam ii4655.CONFIG_DATA = 16'h9999;
      defparam ii4655.PLACE_LOCATION = "NONE";
      defparam ii4655.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4656 ( .DX(nn4656), .F0(yEnd[10]), .F1(\inputctrl1_yAddress__reg[10]|Q_net ), .F2(dummy_abc_3443_), .F3(dummy_abc_3444_) );
      defparam ii4656.CONFIG_DATA = 16'h9999;
      defparam ii4656.PLACE_LOCATION = "NONE";
      defparam ii4656.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4657 ( .DX(nn4657), .F0(dummy_abc_3445_), .F1(dummy_abc_3446_), .F2(dummy_abc_3447_), .F3(dummy_abc_3448_) );
      defparam ii4657.CONFIG_DATA = 16'hFFFF;
      defparam ii4657.PLACE_LOCATION = "NONE";
      defparam ii4657.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_290_ ( 
        .CA( {a_acc_en_cal1_u137_mac, yEnd[10], yEnd[9], yEnd[8], yEnd[7], 
              yEnd[6], yEnd[5], yEnd[4], yEnd[3], yEnd[2], yEnd[1], yEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_118_ ), 
        .DX( {nn4657, nn4656, nn4655, nn4654, nn4653, nn4652, nn4651, nn4650, 
              nn4649, nn4648, nn4647, nn4646} ), 
        .SUM( {\inputctrl1_u43_XORCI_11|SUM_net , dummy_119_, dummy_120_, 
              dummy_121_, dummy_122_, dummy_123_, dummy_124_, dummy_125_, dummy_126_, 
              dummy_127_, dummy_128_, dummy_129_} )
      );
    CS_LUT4_PRIM ii4672 ( .DX(nn4672), .F0(xBgn[0]), .F1(\inputctrl1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_3449_), .F3(dummy_abc_3450_) );
      defparam ii4672.CONFIG_DATA = 16'h9999;
      defparam ii4672.PLACE_LOCATION = "NONE";
      defparam ii4672.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4673 ( .DX(nn4673), .F0(xBgn[1]), .F1(\inputctrl1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_3451_), .F3(dummy_abc_3452_) );
      defparam ii4673.CONFIG_DATA = 16'h9999;
      defparam ii4673.PLACE_LOCATION = "NONE";
      defparam ii4673.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4674 ( .DX(nn4674), .F0(xBgn[2]), .F1(\inputctrl1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_3453_), .F3(dummy_abc_3454_) );
      defparam ii4674.CONFIG_DATA = 16'h9999;
      defparam ii4674.PLACE_LOCATION = "NONE";
      defparam ii4674.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4675 ( .DX(nn4675), .F0(xBgn[3]), .F1(\inputctrl1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_3455_), .F3(dummy_abc_3456_) );
      defparam ii4675.CONFIG_DATA = 16'h9999;
      defparam ii4675.PLACE_LOCATION = "NONE";
      defparam ii4675.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4676 ( .DX(nn4676), .F0(xBgn[4]), .F1(\inputctrl1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_3457_), .F3(dummy_abc_3458_) );
      defparam ii4676.CONFIG_DATA = 16'h9999;
      defparam ii4676.PLACE_LOCATION = "NONE";
      defparam ii4676.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4677 ( .DX(nn4677), .F0(xBgn[5]), .F1(\inputctrl1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_3459_), .F3(dummy_abc_3460_) );
      defparam ii4677.CONFIG_DATA = 16'h9999;
      defparam ii4677.PLACE_LOCATION = "NONE";
      defparam ii4677.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4678 ( .DX(nn4678), .F0(xBgn[6]), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_3461_), .F3(dummy_abc_3462_) );
      defparam ii4678.CONFIG_DATA = 16'h9999;
      defparam ii4678.PLACE_LOCATION = "NONE";
      defparam ii4678.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4679 ( .DX(nn4679), .F0(xBgn[7]), .F1(\inputctrl1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_3463_), .F3(dummy_abc_3464_) );
      defparam ii4679.CONFIG_DATA = 16'h9999;
      defparam ii4679.PLACE_LOCATION = "NONE";
      defparam ii4679.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4680 ( .DX(nn4680), .F0(xBgn[8]), .F1(\inputctrl1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_3465_), .F3(dummy_abc_3466_) );
      defparam ii4680.CONFIG_DATA = 16'h9999;
      defparam ii4680.PLACE_LOCATION = "NONE";
      defparam ii4680.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4681 ( .DX(nn4681), .F0(xBgn[9]), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_3467_), .F3(dummy_abc_3468_) );
      defparam ii4681.CONFIG_DATA = 16'h9999;
      defparam ii4681.PLACE_LOCATION = "NONE";
      defparam ii4681.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4682 ( .DX(nn4682), .F0(xBgn[10]), .F1(\inputctrl1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_3469_), .F3(dummy_abc_3470_) );
      defparam ii4682.CONFIG_DATA = 16'h9999;
      defparam ii4682.PLACE_LOCATION = "NONE";
      defparam ii4682.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4683 ( .DX(nn4683), .F0(dummy_abc_3471_), .F1(dummy_abc_3472_), .F2(dummy_abc_3473_), .F3(dummy_abc_3474_) );
      defparam ii4683.CONFIG_DATA = 16'hFFFF;
      defparam ii4683.PLACE_LOCATION = "NONE";
      defparam ii4683.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_287_ ( 
        .CA( {a_acc_en_cal1_u137_mac, \inputctrl1_xAddress__reg[10]|Q_net , 
              \inputctrl1_xAddress__reg[9]|Q_net , \inputctrl1_xAddress__reg[8]|Q_net , 
              \inputctrl1_xAddress__reg[7]|Q_net , \inputctrl1_xAddress__reg[6]|Q_net , 
              \inputctrl1_xAddress__reg[5]|Q_net , \inputctrl1_xAddress__reg[4]|Q_net , 
              \inputctrl1_xAddress__reg[3]|Q_net , \inputctrl1_xAddress__reg[2]|Q_net , 
              \inputctrl1_xAddress__reg[1]|Q_net , \inputctrl1_xAddress__reg[0]|Q_net } ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_79_ ), 
        .DX( {nn4683, nn4682, nn4681, nn4680, nn4679, nn4678, nn4677, nn4676, 
              nn4675, nn4674, nn4673, nn4672} ), 
        .SUM( {\inputctrl1_u37_XORCI_11|SUM_net , dummy_80_, dummy_81_, dummy_82_, 
              dummy_83_, dummy_84_, dummy_85_, dummy_86_, dummy_87_, dummy_88_, 
              dummy_89_, dummy_90_} )
      );
    CS_LUT4_PRIM ii4698 ( .DX(nn4698), .F0(xEnd[0]), .F1(\inputctrl1_xAddress__reg[0]|Q_net ), .F2(dummy_abc_3475_), .F3(dummy_abc_3476_) );
      defparam ii4698.CONFIG_DATA = 16'h9999;
      defparam ii4698.PLACE_LOCATION = "NONE";
      defparam ii4698.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4699 ( .DX(nn4699), .F0(xEnd[1]), .F1(\inputctrl1_xAddress__reg[1]|Q_net ), .F2(dummy_abc_3477_), .F3(dummy_abc_3478_) );
      defparam ii4699.CONFIG_DATA = 16'h9999;
      defparam ii4699.PLACE_LOCATION = "NONE";
      defparam ii4699.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4700 ( .DX(nn4700), .F0(xEnd[2]), .F1(\inputctrl1_xAddress__reg[2]|Q_net ), .F2(dummy_abc_3479_), .F3(dummy_abc_3480_) );
      defparam ii4700.CONFIG_DATA = 16'h9999;
      defparam ii4700.PLACE_LOCATION = "NONE";
      defparam ii4700.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4701 ( .DX(nn4701), .F0(xEnd[3]), .F1(\inputctrl1_xAddress__reg[3]|Q_net ), .F2(dummy_abc_3481_), .F3(dummy_abc_3482_) );
      defparam ii4701.CONFIG_DATA = 16'h9999;
      defparam ii4701.PLACE_LOCATION = "NONE";
      defparam ii4701.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4702 ( .DX(nn4702), .F0(xEnd[4]), .F1(\inputctrl1_xAddress__reg[4]|Q_net ), .F2(dummy_abc_3483_), .F3(dummy_abc_3484_) );
      defparam ii4702.CONFIG_DATA = 16'h9999;
      defparam ii4702.PLACE_LOCATION = "NONE";
      defparam ii4702.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4703 ( .DX(nn4703), .F0(xEnd[5]), .F1(\inputctrl1_xAddress__reg[5]|Q_net ), .F2(dummy_abc_3485_), .F3(dummy_abc_3486_) );
      defparam ii4703.CONFIG_DATA = 16'h9999;
      defparam ii4703.PLACE_LOCATION = "NONE";
      defparam ii4703.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4704 ( .DX(nn4704), .F0(xEnd[6]), .F1(\inputctrl1_xAddress__reg[6]|Q_net ), .F2(dummy_abc_3487_), .F3(dummy_abc_3488_) );
      defparam ii4704.CONFIG_DATA = 16'h9999;
      defparam ii4704.PLACE_LOCATION = "NONE";
      defparam ii4704.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4705 ( .DX(nn4705), .F0(xEnd[7]), .F1(\inputctrl1_xAddress__reg[7]|Q_net ), .F2(dummy_abc_3489_), .F3(dummy_abc_3490_) );
      defparam ii4705.CONFIG_DATA = 16'h9999;
      defparam ii4705.PLACE_LOCATION = "NONE";
      defparam ii4705.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4706 ( .DX(nn4706), .F0(xEnd[8]), .F1(\inputctrl1_xAddress__reg[8]|Q_net ), .F2(dummy_abc_3491_), .F3(dummy_abc_3492_) );
      defparam ii4706.CONFIG_DATA = 16'h9999;
      defparam ii4706.PLACE_LOCATION = "NONE";
      defparam ii4706.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4707 ( .DX(nn4707), .F0(xEnd[9]), .F1(\inputctrl1_xAddress__reg[9]|Q_net ), .F2(dummy_abc_3493_), .F3(dummy_abc_3494_) );
      defparam ii4707.CONFIG_DATA = 16'h9999;
      defparam ii4707.PLACE_LOCATION = "NONE";
      defparam ii4707.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4708 ( .DX(nn4708), .F0(xEnd[10]), .F1(\inputctrl1_xAddress__reg[10]|Q_net ), .F2(dummy_abc_3495_), .F3(dummy_abc_3496_) );
      defparam ii4708.CONFIG_DATA = 16'h9999;
      defparam ii4708.PLACE_LOCATION = "NONE";
      defparam ii4708.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4709 ( .DX(nn4709), .F0(dummy_abc_3497_), .F1(dummy_abc_3498_), .F2(dummy_abc_3499_), .F3(dummy_abc_3500_) );
      defparam ii4709.CONFIG_DATA = 16'hFFFF;
      defparam ii4709.PLACE_LOCATION = "NONE";
      defparam ii4709.PCK_LOCATION = "NONE";
    scaler_ipc_adder_12 carry_12_289_ ( 
        .CA( {a_acc_en_cal1_u137_mac, xEnd[10], xEnd[9], xEnd[8], xEnd[7], 
              xEnd[6], xEnd[5], xEnd[4], xEnd[3], xEnd[2], xEnd[1], xEnd[0]} ), 
        .CI( a_dinxy_cen_cal1_u137_mac ), 
        .CO( dummy_105_ ), 
        .DX( {nn4709, nn4708, nn4707, nn4706, nn4705, nn4704, nn4703, nn4702, 
              nn4701, nn4700, nn4699, nn4698} ), 
        .SUM( {\inputctrl1_u41_XORCI_11|SUM_net , dummy_106_, dummy_107_, 
              dummy_108_, dummy_109_, dummy_110_, dummy_111_, dummy_112_, dummy_113_, 
              dummy_114_, dummy_115_, dummy_116_} )
      );
    CS_LUT4_PRIM ii4724 ( .DX(nn4724), .F0(dInEn), .F1(dummy_118_), .F2(dummy_79_), .F3(dummy_105_) );
      defparam ii4724.CONFIG_DATA = 16'h8000;
      defparam ii4724.PLACE_LOCATION = "NONE";
      defparam ii4724.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4725 ( .DX(nn4725), .F0(\inputctrl1_yPreEn__reg|Q_net ), .F1(dummy_92_), .F2(nn4645), .F3(nn4724) );
      defparam ii4725.CONFIG_DATA = 16'hC800;
      defparam ii4725.PLACE_LOCATION = "NONE";
      defparam ii4725.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4726 ( .DX(nn4726), .F0(\inputctrl1_xPreEn__reg|Q_net ), .F1(nn4612), .F2(nn4725), .F3(dummy_abc_3501_) );
      defparam ii4726.CONFIG_DATA = 16'hE0E0;
      defparam ii4726.PLACE_LOCATION = "NONE";
      defparam ii4726.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4727 ( .DX(nn4727), .F0(iHsyn), .F1(iVsyn), .F2(nn4726), .F3(dummy_abc_3502_) );
      defparam ii4727.CONFIG_DATA = 16'hFEFE;
      defparam ii4727.PLACE_LOCATION = "NONE";
      defparam ii4727.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4728 ( .DX(nn4728), .F0(dIn[10]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3503_) );
      defparam ii4728.CONFIG_DATA = 16'h0202;
      defparam ii4728.PLACE_LOCATION = "NONE";
      defparam ii4728.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4729 ( .DX(nn4729), .F0(dIn[11]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3504_) );
      defparam ii4729.CONFIG_DATA = 16'h0202;
      defparam ii4729.PLACE_LOCATION = "NONE";
      defparam ii4729.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4730 ( .DX(nn4730), .F0(dIn[12]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3505_) );
      defparam ii4730.CONFIG_DATA = 16'h0202;
      defparam ii4730.PLACE_LOCATION = "NONE";
      defparam ii4730.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4731 ( .DX(nn4731), .F0(dIn[13]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3506_) );
      defparam ii4731.CONFIG_DATA = 16'h0202;
      defparam ii4731.PLACE_LOCATION = "NONE";
      defparam ii4731.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4732 ( .DX(nn4732), .F0(dIn[14]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3507_) );
      defparam ii4732.CONFIG_DATA = 16'h0202;
      defparam ii4732.PLACE_LOCATION = "NONE";
      defparam ii4732.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4733 ( .DX(nn4733), .F0(dIn[15]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3508_) );
      defparam ii4733.CONFIG_DATA = 16'h0202;
      defparam ii4733.PLACE_LOCATION = "NONE";
      defparam ii4733.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4734 ( .DX(nn4734), .F0(dIn[16]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3509_) );
      defparam ii4734.CONFIG_DATA = 16'h0202;
      defparam ii4734.PLACE_LOCATION = "NONE";
      defparam ii4734.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4735 ( .DX(nn4735), .F0(dIn[17]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3510_) );
      defparam ii4735.CONFIG_DATA = 16'h0202;
      defparam ii4735.PLACE_LOCATION = "NONE";
      defparam ii4735.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4736 ( .DX(nn4736), .F0(dIn[18]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3511_) );
      defparam ii4736.CONFIG_DATA = 16'h0202;
      defparam ii4736.PLACE_LOCATION = "NONE";
      defparam ii4736.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4737 ( .DX(nn4737), .F0(dIn[19]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3512_) );
      defparam ii4737.CONFIG_DATA = 16'h0202;
      defparam ii4737.PLACE_LOCATION = "NONE";
      defparam ii4737.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4738 ( .DX(nn4738), .F0(dIn[1]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3513_) );
      defparam ii4738.CONFIG_DATA = 16'h0202;
      defparam ii4738.PLACE_LOCATION = "NONE";
      defparam ii4738.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4739 ( .DX(nn4739), .F0(dIn[20]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3514_) );
      defparam ii4739.CONFIG_DATA = 16'h0202;
      defparam ii4739.PLACE_LOCATION = "NONE";
      defparam ii4739.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4740 ( .DX(nn4740), .F0(dIn[21]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3515_) );
      defparam ii4740.CONFIG_DATA = 16'h0202;
      defparam ii4740.PLACE_LOCATION = "NONE";
      defparam ii4740.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4741 ( .DX(nn4741), .F0(dIn[22]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3516_) );
      defparam ii4741.CONFIG_DATA = 16'h0202;
      defparam ii4741.PLACE_LOCATION = "NONE";
      defparam ii4741.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4742 ( .DX(nn4742), .F0(dIn[23]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3517_) );
      defparam ii4742.CONFIG_DATA = 16'h0202;
      defparam ii4742.PLACE_LOCATION = "NONE";
      defparam ii4742.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4743 ( .DX(nn4743), .F0(dIn[2]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3518_) );
      defparam ii4743.CONFIG_DATA = 16'h0202;
      defparam ii4743.PLACE_LOCATION = "NONE";
      defparam ii4743.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4744 ( .DX(nn4744), .F0(dIn[3]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3519_) );
      defparam ii4744.CONFIG_DATA = 16'h0202;
      defparam ii4744.PLACE_LOCATION = "NONE";
      defparam ii4744.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4745 ( .DX(nn4745), .F0(dIn[4]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3520_) );
      defparam ii4745.CONFIG_DATA = 16'h0202;
      defparam ii4745.PLACE_LOCATION = "NONE";
      defparam ii4745.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4746 ( .DX(nn4746), .F0(dIn[5]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3521_) );
      defparam ii4746.CONFIG_DATA = 16'h0202;
      defparam ii4746.PLACE_LOCATION = "NONE";
      defparam ii4746.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4747 ( .DX(nn4747), .F0(dIn[6]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3522_) );
      defparam ii4747.CONFIG_DATA = 16'h0202;
      defparam ii4747.PLACE_LOCATION = "NONE";
      defparam ii4747.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4748 ( .DX(nn4748), .F0(dIn[7]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3523_) );
      defparam ii4748.CONFIG_DATA = 16'h0202;
      defparam ii4748.PLACE_LOCATION = "NONE";
      defparam ii4748.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4749 ( .DX(nn4749), .F0(dIn[8]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3524_) );
      defparam ii4749.CONFIG_DATA = 16'h0202;
      defparam ii4749.PLACE_LOCATION = "NONE";
      defparam ii4749.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4750 ( .DX(nn4750), .F0(dIn[9]), .F1(iHsyn), .F2(iVsyn), .F3(dummy_abc_3525_) );
      defparam ii4750.CONFIG_DATA = 16'h0202;
      defparam ii4750.PLACE_LOCATION = "NONE";
      defparam ii4750.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4751 ( .DX(nn4751), .F0(iHsyn), .F1(\inputctrl1_yPreEn__reg|Q_net ), .F2(nn4645), .F3(dummy_abc_3526_) );
      defparam ii4751.CONFIG_DATA = 16'hA8A8;
      defparam ii4751.PLACE_LOCATION = "NONE";
      defparam ii4751.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4752 ( .DX(nn4752), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F3(dummy_abc_3527_) );
      defparam ii4752.CONFIG_DATA = 16'hEFEF;
      defparam ii4752.PLACE_LOCATION = "NONE";
      defparam ii4752.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4753 ( .DX(nn4753), .F0(\inputctrl1_ramWrtAddr__reg[0]|Q_net ), .F1(dummy_abc_3528_), .F2(dummy_abc_3529_), .F3(dummy_abc_3530_) );
      defparam ii4753.CONFIG_DATA = 16'h5555;
      defparam ii4753.PLACE_LOCATION = "NONE";
      defparam ii4753.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4754 ( .DX(nn4754), .F0(\inputctrl1_ramWrtAddr__reg[1]|Q_net ), .F1(dummy_abc_3531_), .F2(dummy_abc_3532_), .F3(dummy_abc_3533_) );
      defparam ii4754.CONFIG_DATA = 16'hAAAA;
      defparam ii4754.PLACE_LOCATION = "NONE";
      defparam ii4754.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4755 ( .DX(nn4755), .F0(\inputctrl1_ramWrtAddr__reg[2]|Q_net ), .F1(dummy_abc_3534_), .F2(dummy_abc_3535_), .F3(dummy_abc_3536_) );
      defparam ii4755.CONFIG_DATA = 16'hAAAA;
      defparam ii4755.PLACE_LOCATION = "NONE";
      defparam ii4755.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4756 ( .DX(nn4756), .F0(\inputctrl1_ramWrtAddr__reg[3]|Q_net ), .F1(dummy_abc_3537_), .F2(dummy_abc_3538_), .F3(dummy_abc_3539_) );
      defparam ii4756.CONFIG_DATA = 16'hAAAA;
      defparam ii4756.PLACE_LOCATION = "NONE";
      defparam ii4756.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4757 ( .DX(nn4757), .F0(\inputctrl1_ramWrtAddr__reg[4]|Q_net ), .F1(dummy_abc_3540_), .F2(dummy_abc_3541_), .F3(dummy_abc_3542_) );
      defparam ii4757.CONFIG_DATA = 16'hAAAA;
      defparam ii4757.PLACE_LOCATION = "NONE";
      defparam ii4757.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4758 ( .DX(nn4758), .F0(\inputctrl1_ramWrtAddr__reg[5]|Q_net ), .F1(dummy_abc_3543_), .F2(dummy_abc_3544_), .F3(dummy_abc_3545_) );
      defparam ii4758.CONFIG_DATA = 16'hAAAA;
      defparam ii4758.PLACE_LOCATION = "NONE";
      defparam ii4758.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4759 ( .DX(nn4759), .F0(\inputctrl1_ramWrtAddr__reg[6]|Q_net ), .F1(dummy_abc_3546_), .F2(dummy_abc_3547_), .F3(dummy_abc_3548_) );
      defparam ii4759.CONFIG_DATA = 16'hAAAA;
      defparam ii4759.PLACE_LOCATION = "NONE";
      defparam ii4759.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4760 ( .DX(nn4760), .F0(\inputctrl1_ramWrtAddr__reg[7]|Q_net ), .F1(dummy_abc_3549_), .F2(dummy_abc_3550_), .F3(dummy_abc_3551_) );
      defparam ii4760.CONFIG_DATA = 16'hAAAA;
      defparam ii4760.PLACE_LOCATION = "NONE";
      defparam ii4760.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4761 ( .DX(nn4761), .F0(\inputctrl1_ramWrtAddr__reg[8]|Q_net ), .F1(dummy_abc_3552_), .F2(dummy_abc_3553_), .F3(dummy_abc_3554_) );
      defparam ii4761.CONFIG_DATA = 16'hAAAA;
      defparam ii4761.PLACE_LOCATION = "NONE";
      defparam ii4761.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4762 ( .DX(nn4762), .F0(\inputctrl1_ramWrtAddr__reg[9]|Q_net ), .F1(dummy_abc_3555_), .F2(dummy_abc_3556_), .F3(dummy_abc_3557_) );
      defparam ii4762.CONFIG_DATA = 16'hAAAA;
      defparam ii4762.PLACE_LOCATION = "NONE";
      defparam ii4762.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4763 ( .DX(nn4763), .F0(\inputctrl1_ramWrtAddr__reg[10]|Q_net ), .F1(dummy_abc_3558_), .F2(dummy_abc_3559_), .F3(dummy_abc_3560_) );
      defparam ii4763.CONFIG_DATA = 16'hAAAA;
      defparam ii4763.PLACE_LOCATION = "NONE";
      defparam ii4763.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_286_ ( 
        .CA( {\inputctrl1_ramWrtAddr__reg[10]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[9]|Q_net , \inputctrl1_ramWrtAddr__reg[8]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[7]|Q_net , \inputctrl1_ramWrtAddr__reg[6]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[5]|Q_net , \inputctrl1_ramWrtAddr__reg[4]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[3]|Q_net , \inputctrl1_ramWrtAddr__reg[2]|Q_net , 
              \inputctrl1_ramWrtAddr__reg[1]|Q_net , \inputctrl1_ramWrtAddr__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_21_ ), 
        .DX( {nn4763, nn4762, nn4761, nn4760, nn4759, nn4758, nn4757, nn4756, 
              nn4755, nn4754, nn4753} ), 
        .SUM( {\inputctrl1_u112_XORCI_10|SUM_net , 
              \inputctrl1_u112_XORCI_9|SUM_net , \inputctrl1_u112_XORCI_8|SUM_net , 
              \inputctrl1_u112_XORCI_7|SUM_net , \inputctrl1_u112_XORCI_6|SUM_net , 
              \inputctrl1_u112_XORCI_5|SUM_net , \inputctrl1_u112_XORCI_4|SUM_net , 
              \inputctrl1_u112_XORCI_3|SUM_net , \inputctrl1_u112_XORCI_2|SUM_net , 
              \inputctrl1_u112_XORCI_1|SUM_net , \inputctrl1_u112_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4777 ( .DX(nn4777), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_10|SUM_net ), .F3(dummy_abc_3561_) );
      defparam ii4777.CONFIG_DATA = 16'hFEFE;
      defparam ii4777.PLACE_LOCATION = "NONE";
      defparam ii4777.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4778 ( .DX(nn4778), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_1|SUM_net ), .F3(dummy_abc_3562_) );
      defparam ii4778.CONFIG_DATA = 16'hFEFE;
      defparam ii4778.PLACE_LOCATION = "NONE";
      defparam ii4778.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4779 ( .DX(nn4779), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_2|SUM_net ), .F3(dummy_abc_3563_) );
      defparam ii4779.CONFIG_DATA = 16'hFEFE;
      defparam ii4779.PLACE_LOCATION = "NONE";
      defparam ii4779.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4780 ( .DX(nn4780), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_3|SUM_net ), .F3(dummy_abc_3564_) );
      defparam ii4780.CONFIG_DATA = 16'hFEFE;
      defparam ii4780.PLACE_LOCATION = "NONE";
      defparam ii4780.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4781 ( .DX(nn4781), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_4|SUM_net ), .F3(dummy_abc_3565_) );
      defparam ii4781.CONFIG_DATA = 16'hFEFE;
      defparam ii4781.PLACE_LOCATION = "NONE";
      defparam ii4781.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4782 ( .DX(nn4782), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_5|SUM_net ), .F3(dummy_abc_3566_) );
      defparam ii4782.CONFIG_DATA = 16'hFEFE;
      defparam ii4782.PLACE_LOCATION = "NONE";
      defparam ii4782.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4783 ( .DX(nn4783), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_6|SUM_net ), .F3(dummy_abc_3567_) );
      defparam ii4783.CONFIG_DATA = 16'hFEFE;
      defparam ii4783.PLACE_LOCATION = "NONE";
      defparam ii4783.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4784 ( .DX(nn4784), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_7|SUM_net ), .F3(dummy_abc_3568_) );
      defparam ii4784.CONFIG_DATA = 16'hFEFE;
      defparam ii4784.PLACE_LOCATION = "NONE";
      defparam ii4784.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4785 ( .DX(nn4785), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_8|SUM_net ), .F3(dummy_abc_3569_) );
      defparam ii4785.CONFIG_DATA = 16'hFEFE;
      defparam ii4785.PLACE_LOCATION = "NONE";
      defparam ii4785.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4786 ( .DX(nn4786), .F0(iHsyn), .F1(iVsyn), .F2(\inputctrl1_u112_XORCI_9|SUM_net ), .F3(dummy_abc_3570_) );
      defparam ii4786.CONFIG_DATA = 16'hFEFE;
      defparam ii4786.PLACE_LOCATION = "NONE";
      defparam ii4786.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4787 ( .DX(nn4787), .F0(iHsyn), .F1(iVsyn), .F2(nn4726), .F3(dummy_abc_3571_) );
      defparam ii4787.CONFIG_DATA = 16'h1010;
      defparam ii4787.PLACE_LOCATION = "NONE";
      defparam ii4787.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4788 ( .DX(nn4788), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_3572_), .F2(dummy_abc_3573_), .F3(dummy_abc_3574_) );
      defparam ii4788.CONFIG_DATA = 16'h5555;
      defparam ii4788.PLACE_LOCATION = "NONE";
      defparam ii4788.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4789 ( .DX(nn4789), .F0(iHsyn), .F1(iVsyn), .F2(rst), .F3(\coefcal1_inEn__reg|Q_net ) );
      defparam ii4789.CONFIG_DATA = 16'hFEF0;
      defparam ii4789.PLACE_LOCATION = "NONE";
      defparam ii4789.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4790 ( .DX(nn4790), .F0(dInEn), .F1(\coefcal1_inEn__reg|Q_net ), .F2(dummy_abc_3575_), .F3(dummy_abc_3576_) );
      defparam ii4790.CONFIG_DATA = 16'h8888;
      defparam ii4790.PLACE_LOCATION = "NONE";
      defparam ii4790.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4791 ( .DX(nn4791), .F0(\inputctrl1_xAddress__reg[0]|Q_net ), .F1(dummy_abc_3577_), .F2(dummy_abc_3578_), .F3(dummy_abc_3579_) );
      defparam ii4791.CONFIG_DATA = 16'h5555;
      defparam ii4791.PLACE_LOCATION = "NONE";
      defparam ii4791.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4792 ( .DX(nn4792), .F0(\inputctrl1_xAddress__reg[1]|Q_net ), .F1(dummy_abc_3580_), .F2(dummy_abc_3581_), .F3(dummy_abc_3582_) );
      defparam ii4792.CONFIG_DATA = 16'hAAAA;
      defparam ii4792.PLACE_LOCATION = "NONE";
      defparam ii4792.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4793 ( .DX(nn4793), .F0(\inputctrl1_xAddress__reg[2]|Q_net ), .F1(dummy_abc_3583_), .F2(dummy_abc_3584_), .F3(dummy_abc_3585_) );
      defparam ii4793.CONFIG_DATA = 16'hAAAA;
      defparam ii4793.PLACE_LOCATION = "NONE";
      defparam ii4793.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4794 ( .DX(nn4794), .F0(\inputctrl1_xAddress__reg[3]|Q_net ), .F1(dummy_abc_3586_), .F2(dummy_abc_3587_), .F3(dummy_abc_3588_) );
      defparam ii4794.CONFIG_DATA = 16'hAAAA;
      defparam ii4794.PLACE_LOCATION = "NONE";
      defparam ii4794.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4795 ( .DX(nn4795), .F0(\inputctrl1_xAddress__reg[4]|Q_net ), .F1(dummy_abc_3589_), .F2(dummy_abc_3590_), .F3(dummy_abc_3591_) );
      defparam ii4795.CONFIG_DATA = 16'hAAAA;
      defparam ii4795.PLACE_LOCATION = "NONE";
      defparam ii4795.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4796 ( .DX(nn4796), .F0(\inputctrl1_xAddress__reg[5]|Q_net ), .F1(dummy_abc_3592_), .F2(dummy_abc_3593_), .F3(dummy_abc_3594_) );
      defparam ii4796.CONFIG_DATA = 16'hAAAA;
      defparam ii4796.PLACE_LOCATION = "NONE";
      defparam ii4796.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4797 ( .DX(nn4797), .F0(\inputctrl1_xAddress__reg[6]|Q_net ), .F1(dummy_abc_3595_), .F2(dummy_abc_3596_), .F3(dummy_abc_3597_) );
      defparam ii4797.CONFIG_DATA = 16'hAAAA;
      defparam ii4797.PLACE_LOCATION = "NONE";
      defparam ii4797.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4798 ( .DX(nn4798), .F0(\inputctrl1_xAddress__reg[7]|Q_net ), .F1(dummy_abc_3598_), .F2(dummy_abc_3599_), .F3(dummy_abc_3600_) );
      defparam ii4798.CONFIG_DATA = 16'hAAAA;
      defparam ii4798.PLACE_LOCATION = "NONE";
      defparam ii4798.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4799 ( .DX(nn4799), .F0(\inputctrl1_xAddress__reg[8]|Q_net ), .F1(dummy_abc_3601_), .F2(dummy_abc_3602_), .F3(dummy_abc_3603_) );
      defparam ii4799.CONFIG_DATA = 16'hAAAA;
      defparam ii4799.PLACE_LOCATION = "NONE";
      defparam ii4799.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4800 ( .DX(nn4800), .F0(\inputctrl1_xAddress__reg[9]|Q_net ), .F1(dummy_abc_3604_), .F2(dummy_abc_3605_), .F3(dummy_abc_3606_) );
      defparam ii4800.CONFIG_DATA = 16'hAAAA;
      defparam ii4800.PLACE_LOCATION = "NONE";
      defparam ii4800.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4801 ( .DX(nn4801), .F0(\inputctrl1_xAddress__reg[10]|Q_net ), .F1(dummy_abc_3607_), .F2(dummy_abc_3608_), .F3(dummy_abc_3609_) );
      defparam ii4801.CONFIG_DATA = 16'hAAAA;
      defparam ii4801.PLACE_LOCATION = "NONE";
      defparam ii4801.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_284_ ( 
        .CA( {\inputctrl1_xAddress__reg[10]|Q_net , 
              \inputctrl1_xAddress__reg[9]|Q_net , \inputctrl1_xAddress__reg[8]|Q_net , 
              \inputctrl1_xAddress__reg[7]|Q_net , \inputctrl1_xAddress__reg[6]|Q_net , 
              \inputctrl1_xAddress__reg[5]|Q_net , \inputctrl1_xAddress__reg[4]|Q_net , 
              \inputctrl1_xAddress__reg[3]|Q_net , \inputctrl1_xAddress__reg[2]|Q_net , 
              \inputctrl1_xAddress__reg[1]|Q_net , \inputctrl1_xAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_19_ ), 
        .DX( {nn4801, nn4800, nn4799, nn4798, nn4797, nn4796, nn4795, nn4794, 
              nn4793, nn4792, nn4791} ), 
        .SUM( {\inputctrl1_u110_XORCI_10|SUM_net , 
              \inputctrl1_u110_XORCI_9|SUM_net , \inputctrl1_u110_XORCI_8|SUM_net , 
              \inputctrl1_u110_XORCI_7|SUM_net , \inputctrl1_u110_XORCI_6|SUM_net , 
              \inputctrl1_u110_XORCI_5|SUM_net , \inputctrl1_u110_XORCI_4|SUM_net , 
              \inputctrl1_u110_XORCI_3|SUM_net , \inputctrl1_u110_XORCI_2|SUM_net , 
              \inputctrl1_u110_XORCI_1|SUM_net , \inputctrl1_u110_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4815 ( .DX(nn4815), .F0(\coefcal1_u61_XORCI_6|SUM_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_79_), .F3(dummy_abc_3610_) );
      defparam ii4815.CONFIG_DATA = 16'hE0E0;
      defparam ii4815.PLACE_LOCATION = "NONE";
      defparam ii4815.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4816 ( .DX(nn4816), .F0(\inputctrl1_xCal__reg[0]|Q_net ), .F1(nn4216), .F2(nn4815), .F3(dummy_abc_3611_) );
      defparam ii4816.CONFIG_DATA = 16'h6A6A;
      defparam ii4816.PLACE_LOCATION = "NONE";
      defparam ii4816.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4817 ( .DX(nn4817), .F0(nn4612), .F1(nn4790), .F2(dummy_abc_3612_), .F3(dummy_abc_3613_) );
      defparam ii4817.CONFIG_DATA = 16'h8888;
      defparam ii4817.PLACE_LOCATION = "NONE";
      defparam ii4817.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4818 ( .DX(nn4818), .F0(\inputctrl1_xCal__reg[0]|Q_net ), .F1(nn4216), .F2(nn4815), .F3(dummy_abc_3614_) );
      defparam ii4818.CONFIG_DATA = 16'h6A6A;
      defparam ii4818.PLACE_LOCATION = "NONE";
      defparam ii4818.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4819 ( .DX(nn4819), .F0(\inputctrl1_xCal__reg[1]|Q_net ), .F1(\coefcal1_u61_XORCI_1|SUM_net ), .F2(nn4815), .F3(dummy_abc_3615_) );
      defparam ii4819.CONFIG_DATA = 16'h6A6A;
      defparam ii4819.PLACE_LOCATION = "NONE";
      defparam ii4819.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4820 ( .DX(nn4820), .F0(\inputctrl1_xCal__reg[2]|Q_net ), .F1(\coefcal1_u61_XORCI_2|SUM_net ), .F2(nn4815), .F3(dummy_abc_3616_) );
      defparam ii4820.CONFIG_DATA = 16'h6A6A;
      defparam ii4820.PLACE_LOCATION = "NONE";
      defparam ii4820.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4821 ( .DX(nn4821), .F0(\inputctrl1_xCal__reg[3]|Q_net ), .F1(\coefcal1_u61_XORCI_3|SUM_net ), .F2(nn4815), .F3(dummy_abc_3617_) );
      defparam ii4821.CONFIG_DATA = 16'h6A6A;
      defparam ii4821.PLACE_LOCATION = "NONE";
      defparam ii4821.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4822 ( .DX(nn4822), .F0(\inputctrl1_xCal__reg[4]|Q_net ), .F1(\coefcal1_u61_XORCI_4|SUM_net ), .F2(nn4815), .F3(dummy_abc_3618_) );
      defparam ii4822.CONFIG_DATA = 16'h6A6A;
      defparam ii4822.PLACE_LOCATION = "NONE";
      defparam ii4822.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4823 ( .DX(nn4823), .F0(\inputctrl1_xCal__reg[5]|Q_net ), .F1(\coefcal1_u61_XORCI_5|SUM_net ), .F2(nn4815), .F3(dummy_abc_3619_) );
      defparam ii4823.CONFIG_DATA = 16'h6A6A;
      defparam ii4823.PLACE_LOCATION = "NONE";
      defparam ii4823.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4824 ( .DX(nn4824), .F0(\inputctrl1_xCal__reg[6]|Q_net ), .F1(\coefcal1_u61_XORCI_6|SUM_net ), .F2(nn4815), .F3(dummy_abc_3620_) );
      defparam ii4824.CONFIG_DATA = 16'h6565;
      defparam ii4824.PLACE_LOCATION = "NONE";
      defparam ii4824.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4825 ( .DX(nn4825), .F0(\inputctrl1_xCal__reg[7]|Q_net ), .F1(\coefcal1_u61_XORCI_7|SUM_net ), .F2(dummy_79_), .F3(dummy_abc_3621_) );
      defparam ii4825.CONFIG_DATA = 16'h6A6A;
      defparam ii4825.PLACE_LOCATION = "NONE";
      defparam ii4825.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4826 ( .DX(nn4826), .F0(\inputctrl1_xCal__reg[8]|Q_net ), .F1(dummy_abc_3622_), .F2(dummy_abc_3623_), .F3(dummy_abc_3624_) );
      defparam ii4826.CONFIG_DATA = 16'hAAAA;
      defparam ii4826.PLACE_LOCATION = "NONE";
      defparam ii4826.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4827 ( .DX(nn4827), .F0(\inputctrl1_xCal__reg[9]|Q_net ), .F1(dummy_abc_3625_), .F2(dummy_abc_3626_), .F3(dummy_abc_3627_) );
      defparam ii4827.CONFIG_DATA = 16'hAAAA;
      defparam ii4827.PLACE_LOCATION = "NONE";
      defparam ii4827.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4828 ( .DX(nn4828), .F0(\inputctrl1_xCal__reg[10]|Q_net ), .F1(dummy_abc_3628_), .F2(dummy_abc_3629_), .F3(dummy_abc_3630_) );
      defparam ii4828.CONFIG_DATA = 16'hAAAA;
      defparam ii4828.PLACE_LOCATION = "NONE";
      defparam ii4828.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4829 ( .DX(nn4829), .F0(\inputctrl1_xCal__reg[11]|Q_net ), .F1(dummy_abc_3631_), .F2(dummy_abc_3632_), .F3(dummy_abc_3633_) );
      defparam ii4829.CONFIG_DATA = 16'hAAAA;
      defparam ii4829.PLACE_LOCATION = "NONE";
      defparam ii4829.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4830 ( .DX(nn4830), .F0(\inputctrl1_xCal__reg[12]|Q_net ), .F1(dummy_abc_3634_), .F2(dummy_abc_3635_), .F3(dummy_abc_3636_) );
      defparam ii4830.CONFIG_DATA = 16'hAAAA;
      defparam ii4830.PLACE_LOCATION = "NONE";
      defparam ii4830.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4831 ( .DX(nn4831), .F0(\inputctrl1_xCal__reg[13]|Q_net ), .F1(dummy_abc_3637_), .F2(dummy_abc_3638_), .F3(dummy_abc_3639_) );
      defparam ii4831.CONFIG_DATA = 16'hAAAA;
      defparam ii4831.PLACE_LOCATION = "NONE";
      defparam ii4831.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4832 ( .DX(nn4832), .F0(\inputctrl1_xCal__reg[14]|Q_net ), .F1(dummy_abc_3640_), .F2(dummy_abc_3641_), .F3(dummy_abc_3642_) );
      defparam ii4832.CONFIG_DATA = 16'hAAAA;
      defparam ii4832.PLACE_LOCATION = "NONE";
      defparam ii4832.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4833 ( .DX(nn4833), .F0(\inputctrl1_xCal__reg[15]|Q_net ), .F1(dummy_abc_3643_), .F2(dummy_abc_3644_), .F3(dummy_abc_3645_) );
      defparam ii4833.CONFIG_DATA = 16'hAAAA;
      defparam ii4833.PLACE_LOCATION = "NONE";
      defparam ii4833.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4834 ( .DX(nn4834), .F0(\inputctrl1_xCal__reg[16]|Q_net ), .F1(dummy_abc_3646_), .F2(dummy_abc_3647_), .F3(dummy_abc_3648_) );
      defparam ii4834.CONFIG_DATA = 16'hAAAA;
      defparam ii4834.PLACE_LOCATION = "NONE";
      defparam ii4834.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_282_ ( 
        .CA( {\inputctrl1_xCal__reg[16]|Q_net , \inputctrl1_xCal__reg[15]|Q_net , 
              \inputctrl1_xCal__reg[14]|Q_net , \inputctrl1_xCal__reg[13]|Q_net , 
              \inputctrl1_xCal__reg[12]|Q_net , \inputctrl1_xCal__reg[11]|Q_net , 
              \inputctrl1_xCal__reg[10]|Q_net , \inputctrl1_xCal__reg[9]|Q_net , 
              \inputctrl1_xCal__reg[8]|Q_net , \inputctrl1_xCal__reg[7]|Q_net , 
              \inputctrl1_xCal__reg[6]|Q_net , \inputctrl1_xCal__reg[5]|Q_net , 
              \inputctrl1_xCal__reg[4]|Q_net , \inputctrl1_xCal__reg[3]|Q_net , 
              \inputctrl1_xCal__reg[2]|Q_net , \inputctrl1_xCal__reg[1]|Q_net , 
              \inputctrl1_xCal__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_201_ ), 
        .DX( {nn4834, nn4833, nn4832, nn4831, nn4830, nn4829, nn4828, nn4827, 
              nn4826, nn4825, nn4824, nn4823, nn4822, nn4821, nn4820, nn4819, 
              nn4818} ), 
        .SUM( {\inputctrl1_u108_XORCI_16|SUM_net , 
              \inputctrl1_u108_XORCI_15|SUM_net , \inputctrl1_u108_XORCI_14|SUM_net , 
              \inputctrl1_u108_XORCI_13|SUM_net , \inputctrl1_u108_XORCI_12|SUM_net , 
              \inputctrl1_u108_XORCI_11|SUM_net , \inputctrl1_u108_XORCI_10|SUM_net , 
              \inputctrl1_u108_XORCI_9|SUM_net , \inputctrl1_u108_XORCI_8|SUM_net , 
              \inputctrl1_u108_XORCI_7|SUM_net , \inputctrl1_u108_XORCI_6|SUM_net , 
              \inputctrl1_u108_XORCI_5|SUM_net , \inputctrl1_u108_XORCI_4|SUM_net , 
              \inputctrl1_u108_XORCI_3|SUM_net , \inputctrl1_u108_XORCI_2|SUM_net , 
              \inputctrl1_u108_XORCI_1|SUM_net , \inputctrl1_u108_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4854 ( .DX(nn4854), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_3649_), .F2(dummy_abc_3650_), .F3(dummy_abc_3651_) );
      defparam ii4854.CONFIG_DATA = 16'h5555;
      defparam ii4854.PLACE_LOCATION = "NONE";
      defparam ii4854.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4855 ( .DX(nn4855), .F0(iVsyn), .F1(rst), .F2(\coefcal1_inEn__reg|Q_net ), .F3(dummy_abc_3652_) );
      defparam ii4855.CONFIG_DATA = 16'hECEC;
      defparam ii4855.PLACE_LOCATION = "NONE";
      defparam ii4855.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4856 ( .DX(nn4856), .F0(\inputctrl1_yAddress__reg[0]|Q_net ), .F1(dummy_abc_3653_), .F2(dummy_abc_3654_), .F3(dummy_abc_3655_) );
      defparam ii4856.CONFIG_DATA = 16'h5555;
      defparam ii4856.PLACE_LOCATION = "NONE";
      defparam ii4856.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4857 ( .DX(nn4857), .F0(\inputctrl1_yAddress__reg[1]|Q_net ), .F1(dummy_abc_3656_), .F2(dummy_abc_3657_), .F3(dummy_abc_3658_) );
      defparam ii4857.CONFIG_DATA = 16'hAAAA;
      defparam ii4857.PLACE_LOCATION = "NONE";
      defparam ii4857.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4858 ( .DX(nn4858), .F0(\inputctrl1_yAddress__reg[2]|Q_net ), .F1(dummy_abc_3659_), .F2(dummy_abc_3660_), .F3(dummy_abc_3661_) );
      defparam ii4858.CONFIG_DATA = 16'hAAAA;
      defparam ii4858.PLACE_LOCATION = "NONE";
      defparam ii4858.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4859 ( .DX(nn4859), .F0(\inputctrl1_yAddress__reg[3]|Q_net ), .F1(dummy_abc_3662_), .F2(dummy_abc_3663_), .F3(dummy_abc_3664_) );
      defparam ii4859.CONFIG_DATA = 16'hAAAA;
      defparam ii4859.PLACE_LOCATION = "NONE";
      defparam ii4859.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4860 ( .DX(nn4860), .F0(\inputctrl1_yAddress__reg[4]|Q_net ), .F1(dummy_abc_3665_), .F2(dummy_abc_3666_), .F3(dummy_abc_3667_) );
      defparam ii4860.CONFIG_DATA = 16'hAAAA;
      defparam ii4860.PLACE_LOCATION = "NONE";
      defparam ii4860.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4861 ( .DX(nn4861), .F0(\inputctrl1_yAddress__reg[5]|Q_net ), .F1(dummy_abc_3668_), .F2(dummy_abc_3669_), .F3(dummy_abc_3670_) );
      defparam ii4861.CONFIG_DATA = 16'hAAAA;
      defparam ii4861.PLACE_LOCATION = "NONE";
      defparam ii4861.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4862 ( .DX(nn4862), .F0(\inputctrl1_yAddress__reg[6]|Q_net ), .F1(dummy_abc_3671_), .F2(dummy_abc_3672_), .F3(dummy_abc_3673_) );
      defparam ii4862.CONFIG_DATA = 16'hAAAA;
      defparam ii4862.PLACE_LOCATION = "NONE";
      defparam ii4862.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4863 ( .DX(nn4863), .F0(\inputctrl1_yAddress__reg[7]|Q_net ), .F1(dummy_abc_3674_), .F2(dummy_abc_3675_), .F3(dummy_abc_3676_) );
      defparam ii4863.CONFIG_DATA = 16'hAAAA;
      defparam ii4863.PLACE_LOCATION = "NONE";
      defparam ii4863.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4864 ( .DX(nn4864), .F0(\inputctrl1_yAddress__reg[8]|Q_net ), .F1(dummy_abc_3677_), .F2(dummy_abc_3678_), .F3(dummy_abc_3679_) );
      defparam ii4864.CONFIG_DATA = 16'hAAAA;
      defparam ii4864.PLACE_LOCATION = "NONE";
      defparam ii4864.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4865 ( .DX(nn4865), .F0(\inputctrl1_yAddress__reg[9]|Q_net ), .F1(dummy_abc_3680_), .F2(dummy_abc_3681_), .F3(dummy_abc_3682_) );
      defparam ii4865.CONFIG_DATA = 16'hAAAA;
      defparam ii4865.PLACE_LOCATION = "NONE";
      defparam ii4865.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4866 ( .DX(nn4866), .F0(\inputctrl1_yAddress__reg[10]|Q_net ), .F1(dummy_abc_3683_), .F2(dummy_abc_3684_), .F3(dummy_abc_3685_) );
      defparam ii4866.CONFIG_DATA = 16'hAAAA;
      defparam ii4866.PLACE_LOCATION = "NONE";
      defparam ii4866.PCK_LOCATION = "NONE";
    scaler_ipc_adder_11 carry_11_285_ ( 
        .CA( {\inputctrl1_yAddress__reg[10]|Q_net , 
              \inputctrl1_yAddress__reg[9]|Q_net , \inputctrl1_yAddress__reg[8]|Q_net , 
              \inputctrl1_yAddress__reg[7]|Q_net , \inputctrl1_yAddress__reg[6]|Q_net , 
              \inputctrl1_yAddress__reg[5]|Q_net , \inputctrl1_yAddress__reg[4]|Q_net , 
              \inputctrl1_yAddress__reg[3]|Q_net , \inputctrl1_yAddress__reg[2]|Q_net , 
              \inputctrl1_yAddress__reg[1]|Q_net , \inputctrl1_yAddress__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_20_ ), 
        .DX( {nn4866, nn4865, nn4864, nn4863, nn4862, nn4861, nn4860, nn4859, 
              nn4858, nn4857, nn4856} ), 
        .SUM( {\inputctrl1_u111_XORCI_10|SUM_net , 
              \inputctrl1_u111_XORCI_9|SUM_net , \inputctrl1_u111_XORCI_8|SUM_net , 
              \inputctrl1_u111_XORCI_7|SUM_net , \inputctrl1_u111_XORCI_6|SUM_net , 
              \inputctrl1_u111_XORCI_5|SUM_net , \inputctrl1_u111_XORCI_4|SUM_net , 
              \inputctrl1_u111_XORCI_3|SUM_net , \inputctrl1_u111_XORCI_2|SUM_net , 
              \inputctrl1_u111_XORCI_1|SUM_net , \inputctrl1_u111_XORCI_0|SUM_net } )
      );
    CS_LUT4_PRIM ii4880 ( .DX(nn4880), .F0(nn2835), .F1(\coefcal1_u62_XORCI_6|SUM_net ), .F2(\coefcal1_u62_XORCI_7|SUM_net ), .F3(dummy_92_) );
      defparam ii4880.CONFIG_DATA = 16'hA800;
      defparam ii4880.PLACE_LOCATION = "NONE";
      defparam ii4880.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4881 ( .DX(nn4881), .F0(\inputctrl1_yCal__reg[0]|Q_net ), .F1(nn4880), .F2(dummy_abc_3686_), .F3(dummy_abc_3687_) );
      defparam ii4881.CONFIG_DATA = 16'h6666;
      defparam ii4881.PLACE_LOCATION = "NONE";
      defparam ii4881.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4882 ( .DX(nn4882), .F0(iHsyn), .F1(nn4645), .F2(dummy_abc_3688_), .F3(dummy_abc_3689_) );
      defparam ii4882.CONFIG_DATA = 16'h8888;
      defparam ii4882.PLACE_LOCATION = "NONE";
      defparam ii4882.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4883 ( .DX(nn4883), .F0(\inputctrl1_yCal__reg[0]|Q_net ), .F1(nn4880), .F2(dummy_abc_3690_), .F3(dummy_abc_3691_) );
      defparam ii4883.CONFIG_DATA = 16'h6666;
      defparam ii4883.PLACE_LOCATION = "NONE";
      defparam ii4883.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4884 ( .DX(nn4884), .F0(\coefcal1_u62_XORCI_6|SUM_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_92_), .F3(dummy_abc_3692_) );
      defparam ii4884.CONFIG_DATA = 16'hE0E0;
      defparam ii4884.PLACE_LOCATION = "NONE";
      defparam ii4884.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4885 ( .DX(nn4885), .F0(\inputctrl1_yCal__reg[1]|Q_net ), .F1(\coefcal1_u62_XORCI_1|SUM_net ), .F2(nn4884), .F3(dummy_abc_3693_) );
      defparam ii4885.CONFIG_DATA = 16'h6A6A;
      defparam ii4885.PLACE_LOCATION = "NONE";
      defparam ii4885.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4886 ( .DX(nn4886), .F0(\inputctrl1_yCal__reg[2]|Q_net ), .F1(\coefcal1_u62_XORCI_2|SUM_net ), .F2(nn4884), .F3(dummy_abc_3694_) );
      defparam ii4886.CONFIG_DATA = 16'h6A6A;
      defparam ii4886.PLACE_LOCATION = "NONE";
      defparam ii4886.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4887 ( .DX(nn4887), .F0(\inputctrl1_yCal__reg[3]|Q_net ), .F1(\coefcal1_u62_XORCI_3|SUM_net ), .F2(nn4884), .F3(dummy_abc_3695_) );
      defparam ii4887.CONFIG_DATA = 16'h6A6A;
      defparam ii4887.PLACE_LOCATION = "NONE";
      defparam ii4887.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4888 ( .DX(nn4888), .F0(\inputctrl1_yCal__reg[4]|Q_net ), .F1(\coefcal1_u62_XORCI_4|SUM_net ), .F2(nn4884), .F3(dummy_abc_3696_) );
      defparam ii4888.CONFIG_DATA = 16'h6A6A;
      defparam ii4888.PLACE_LOCATION = "NONE";
      defparam ii4888.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4889 ( .DX(nn4889), .F0(\inputctrl1_yCal__reg[5]|Q_net ), .F1(\coefcal1_u62_XORCI_5|SUM_net ), .F2(nn4884), .F3(dummy_abc_3697_) );
      defparam ii4889.CONFIG_DATA = 16'h6A6A;
      defparam ii4889.PLACE_LOCATION = "NONE";
      defparam ii4889.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4890 ( .DX(nn4890), .F0(\inputctrl1_yCal__reg[6]|Q_net ), .F1(\coefcal1_u62_XORCI_6|SUM_net ), .F2(nn4884), .F3(dummy_abc_3698_) );
      defparam ii4890.CONFIG_DATA = 16'h6565;
      defparam ii4890.PLACE_LOCATION = "NONE";
      defparam ii4890.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4891 ( .DX(nn4891), .F0(\inputctrl1_yCal__reg[7]|Q_net ), .F1(\coefcal1_u62_XORCI_7|SUM_net ), .F2(dummy_92_), .F3(dummy_abc_3699_) );
      defparam ii4891.CONFIG_DATA = 16'h6A6A;
      defparam ii4891.PLACE_LOCATION = "NONE";
      defparam ii4891.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4892 ( .DX(nn4892), .F0(\inputctrl1_yCal__reg[8]|Q_net ), .F1(dummy_abc_3700_), .F2(dummy_abc_3701_), .F3(dummy_abc_3702_) );
      defparam ii4892.CONFIG_DATA = 16'hAAAA;
      defparam ii4892.PLACE_LOCATION = "NONE";
      defparam ii4892.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4893 ( .DX(nn4893), .F0(\inputctrl1_yCal__reg[9]|Q_net ), .F1(dummy_abc_3703_), .F2(dummy_abc_3704_), .F3(dummy_abc_3705_) );
      defparam ii4893.CONFIG_DATA = 16'hAAAA;
      defparam ii4893.PLACE_LOCATION = "NONE";
      defparam ii4893.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4894 ( .DX(nn4894), .F0(\inputctrl1_yCal__reg[10]|Q_net ), .F1(dummy_abc_3706_), .F2(dummy_abc_3707_), .F3(dummy_abc_3708_) );
      defparam ii4894.CONFIG_DATA = 16'hAAAA;
      defparam ii4894.PLACE_LOCATION = "NONE";
      defparam ii4894.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4895 ( .DX(nn4895), .F0(\inputctrl1_yCal__reg[11]|Q_net ), .F1(dummy_abc_3709_), .F2(dummy_abc_3710_), .F3(dummy_abc_3711_) );
      defparam ii4895.CONFIG_DATA = 16'hAAAA;
      defparam ii4895.PLACE_LOCATION = "NONE";
      defparam ii4895.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4896 ( .DX(nn4896), .F0(\inputctrl1_yCal__reg[12]|Q_net ), .F1(dummy_abc_3712_), .F2(dummy_abc_3713_), .F3(dummy_abc_3714_) );
      defparam ii4896.CONFIG_DATA = 16'hAAAA;
      defparam ii4896.PLACE_LOCATION = "NONE";
      defparam ii4896.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4897 ( .DX(nn4897), .F0(\inputctrl1_yCal__reg[13]|Q_net ), .F1(dummy_abc_3715_), .F2(dummy_abc_3716_), .F3(dummy_abc_3717_) );
      defparam ii4897.CONFIG_DATA = 16'hAAAA;
      defparam ii4897.PLACE_LOCATION = "NONE";
      defparam ii4897.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4898 ( .DX(nn4898), .F0(\inputctrl1_yCal__reg[14]|Q_net ), .F1(dummy_abc_3718_), .F2(dummy_abc_3719_), .F3(dummy_abc_3720_) );
      defparam ii4898.CONFIG_DATA = 16'hAAAA;
      defparam ii4898.PLACE_LOCATION = "NONE";
      defparam ii4898.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4899 ( .DX(nn4899), .F0(\inputctrl1_yCal__reg[15]|Q_net ), .F1(dummy_abc_3721_), .F2(dummy_abc_3722_), .F3(dummy_abc_3723_) );
      defparam ii4899.CONFIG_DATA = 16'hAAAA;
      defparam ii4899.PLACE_LOCATION = "NONE";
      defparam ii4899.PCK_LOCATION = "NONE";
    CS_LUT4_PRIM ii4900 ( .DX(nn4900), .F0(\inputctrl1_yCal__reg[16]|Q_net ), .F1(dummy_abc_3724_), .F2(dummy_abc_3725_), .F3(dummy_abc_3726_) );
      defparam ii4900.CONFIG_DATA = 16'hAAAA;
      defparam ii4900.PLACE_LOCATION = "NONE";
      defparam ii4900.PCK_LOCATION = "NONE";
    scaler_ipc_adder_17 carry_17_283_ ( 
        .CA( {\inputctrl1_yCal__reg[16]|Q_net , \inputctrl1_yCal__reg[15]|Q_net , 
              \inputctrl1_yCal__reg[14]|Q_net , \inputctrl1_yCal__reg[13]|Q_net , 
              \inputctrl1_yCal__reg[12]|Q_net , \inputctrl1_yCal__reg[11]|Q_net , 
              \inputctrl1_yCal__reg[10]|Q_net , \inputctrl1_yCal__reg[9]|Q_net , 
              \inputctrl1_yCal__reg[8]|Q_net , \inputctrl1_yCal__reg[7]|Q_net , 
              \inputctrl1_yCal__reg[6]|Q_net , \inputctrl1_yCal__reg[5]|Q_net , 
              \inputctrl1_yCal__reg[4]|Q_net , \inputctrl1_yCal__reg[3]|Q_net , 
              \inputctrl1_yCal__reg[2]|Q_net , \inputctrl1_yCal__reg[1]|Q_net , 
              \inputctrl1_yCal__reg[0]|Q_net } ), 
        .CI( a_acc_en_cal1_u137_mac ), 
        .CO( dummy_202_ ), 
        .DX( {nn4900, nn4899, nn4898, nn4897, nn4896, nn4895, nn4894, nn4893, 
              nn4892, nn4891, nn4890, nn4889, nn4888, nn4887, nn4886, nn4885, 
              nn4883} ), 
        .SUM( {\inputctrl1_u109_XORCI_16|SUM_net , 
              \inputctrl1_u109_XORCI_15|SUM_net , \inputctrl1_u109_XORCI_14|SUM_net , 
              \inputctrl1_u109_XORCI_13|SUM_net , \inputctrl1_u109_XORCI_12|SUM_net , 
              \inputctrl1_u109_XORCI_11|SUM_net , \inputctrl1_u109_XORCI_10|SUM_net , 
              \inputctrl1_u109_XORCI_9|SUM_net , \inputctrl1_u109_XORCI_8|SUM_net , 
              \inputctrl1_u109_XORCI_7|SUM_net , \inputctrl1_u109_XORCI_6|SUM_net , 
              \inputctrl1_u109_XORCI_5|SUM_net , \inputctrl1_u109_XORCI_4|SUM_net , 
              \inputctrl1_u109_XORCI_3|SUM_net , \inputctrl1_u109_XORCI_2|SUM_net , 
              \inputctrl1_u109_XORCI_1|SUM_net , \inputctrl1_u109_XORCI_0|SUM_net } )
      );
    CS_REGA_PRIM cal1_HS__reg ( .CLK( clkb ), .D( nn1517 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( HS_2079_net ) );
      defparam cal1_HS__reg.INIT = 0;
      defparam cal1_HS__reg.PLACE_LOCATION = "NONE";
      defparam cal1_HS__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_VSNormal__reg ( .CLK( clkb ), .D( nn1519 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \cal1_VSNormal__reg|Q_net  ) );
      defparam cal1_VSNormal__reg.INIT = 0;
      defparam cal1_VSNormal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_VSNormal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_enforceJmp__reg ( .CLK( clkb ), .D( a_acc_en_cal1_u137_mac ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \cal1_enforceJmp__reg|Q_net  ) );
      defparam cal1_enforceJmp__reg.INIT = 0;
      defparam cal1_enforceJmp__reg.PLACE_LOCATION = "NONE";
      defparam cal1_enforceJmp__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_jmp1Normal__reg ( .CLK( clkb ), .D( nn2901 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \cal1_jmp1Normal__reg|Q_net  ) );
      defparam cal1_jmp1Normal__reg.INIT = 0;
      defparam cal1_jmp1Normal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_jmp1Normal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM cal1_jmp2Normal__reg ( .CLK( clkb ), .D( nn2902 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \cal1_jmp2Normal__reg|Q_net  ) );
      defparam cal1_jmp2Normal__reg.INIT = 0;
      defparam cal1_jmp2Normal__reg.PLACE_LOCATION = "NONE";
      defparam cal1_jmp2Normal__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[0]  ( .CLK( clkb ), .D( nn4282 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[0]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[0] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[10]  ( .CLK( clkb ), .D( nn4309 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[10]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[10] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[1]  ( .CLK( clkb ), .D( nn4310 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[1]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[1] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[2]  ( .CLK( clkb ), .D( nn4311 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[2]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[2] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[3]  ( .CLK( clkb ), .D( nn4312 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[3]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[3] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[4]  ( .CLK( clkb ), .D( nn4313 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[4]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[4] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[5]  ( .CLK( clkb ), .D( nn4314 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[5]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[5] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[6]  ( .CLK( clkb ), .D( nn4315 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[6]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[6] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[7]  ( .CLK( clkb ), .D( nn4316 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[7]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[7] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[8]  ( .CLK( clkb ), .D( nn4317 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[8]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[8] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_ramRdAddr__reg[9]  ( .CLK( clkb ), .D( nn4318 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4284 ), .Q( \cal1_ramRdAddr__reg[9]|Q_net  ) );
      defparam \cal1_ramRdAddr__reg[9] .INIT = 0;
      defparam \cal1_ramRdAddr__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_ramRdAddr__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[0]  ( .CLK( clkb ), .D( \cal1_u__reg[0]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[0]|Q_net  ) );
      defparam \cal1_uPreF__reg[0] .INIT = 0;
      defparam \cal1_uPreF__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[1]  ( .CLK( clkb ), .D( \cal1_u__reg[1]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[1]|Q_net  ) );
      defparam \cal1_uPreF__reg[1] .INIT = 0;
      defparam \cal1_uPreF__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[2]  ( .CLK( clkb ), .D( \cal1_u__reg[2]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[2]|Q_net  ) );
      defparam \cal1_uPreF__reg[2] .INIT = 0;
      defparam \cal1_uPreF__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[3]  ( .CLK( clkb ), .D( \cal1_u__reg[3]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[3]|Q_net  ) );
      defparam \cal1_uPreF__reg[3] .INIT = 0;
      defparam \cal1_uPreF__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[4]  ( .CLK( clkb ), .D( \cal1_u__reg[4]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[4]|Q_net  ) );
      defparam \cal1_uPreF__reg[4] .INIT = 0;
      defparam \cal1_uPreF__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_uPreF__reg[5]  ( .CLK( clkb ), .D( \cal1_u__reg[5]|Q_net  ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_uPreF__reg[5]|Q_net  ) );
      defparam \cal1_uPreF__reg[5] .INIT = 0;
      defparam \cal1_uPreF__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_uPreF__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[0]  ( .CLK( clkb ), .D( nn4320 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[0]|Q_net  ) );
      defparam \cal1_u__reg[0] .INIT = 0;
      defparam \cal1_u__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[10]  ( .CLK( clkb ), .D( nn4321 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[10]|Q_net  ) );
      defparam \cal1_u__reg[10] .INIT = 0;
      defparam \cal1_u__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[11]  ( .CLK( clkb ), .D( nn4322 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[11]|Q_net  ) );
      defparam \cal1_u__reg[11] .INIT = 0;
      defparam \cal1_u__reg[11] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[12]  ( .CLK( clkb ), .D( nn4323 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[12]|Q_net  ) );
      defparam \cal1_u__reg[12] .INIT = 0;
      defparam \cal1_u__reg[12] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[13]  ( .CLK( clkb ), .D( nn4324 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[13]|Q_net  ) );
      defparam \cal1_u__reg[13] .INIT = 0;
      defparam \cal1_u__reg[13] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[14]  ( .CLK( clkb ), .D( nn4325 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[14]|Q_net  ) );
      defparam \cal1_u__reg[14] .INIT = 0;
      defparam \cal1_u__reg[14] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[15]  ( .CLK( clkb ), .D( nn4326 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[15]|Q_net  ) );
      defparam \cal1_u__reg[15] .INIT = 0;
      defparam \cal1_u__reg[15] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[16]  ( .CLK( clkb ), .D( nn4327 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[16]|Q_net  ) );
      defparam \cal1_u__reg[16] .INIT = 0;
      defparam \cal1_u__reg[16] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[1]  ( .CLK( clkb ), .D( nn4328 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[1]|Q_net  ) );
      defparam \cal1_u__reg[1] .INIT = 0;
      defparam \cal1_u__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[2]  ( .CLK( clkb ), .D( nn4329 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[2]|Q_net  ) );
      defparam \cal1_u__reg[2] .INIT = 0;
      defparam \cal1_u__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[3]  ( .CLK( clkb ), .D( nn4330 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[3]|Q_net  ) );
      defparam \cal1_u__reg[3] .INIT = 0;
      defparam \cal1_u__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[4]  ( .CLK( clkb ), .D( nn4331 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[4]|Q_net  ) );
      defparam \cal1_u__reg[4] .INIT = 0;
      defparam \cal1_u__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[5]  ( .CLK( clkb ), .D( nn4332 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[5]|Q_net  ) );
      defparam \cal1_u__reg[5] .INIT = 0;
      defparam \cal1_u__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[6]  ( .CLK( clkb ), .D( nn4333 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[6]|Q_net  ) );
      defparam \cal1_u__reg[6] .INIT = 0;
      defparam \cal1_u__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[7]  ( .CLK( clkb ), .D( nn4334 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[7]|Q_net  ) );
      defparam \cal1_u__reg[7] .INIT = 0;
      defparam \cal1_u__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[8]  ( .CLK( clkb ), .D( nn4335 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[8]|Q_net  ) );
      defparam \cal1_u__reg[8] .INIT = 0;
      defparam \cal1_u__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_u__reg[9]  ( .CLK( clkb ), .D( nn4336 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_u__reg[9]|Q_net  ) );
      defparam \cal1_u__reg[9] .INIT = 0;
      defparam \cal1_u__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_u__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[0]  ( .CLK( clkb ), .D( nn4338 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[0]|Q_net  ) );
      defparam \cal1_v__reg[0] .INIT = 0;
      defparam \cal1_v__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[10]  ( .CLK( clkb ), .D( nn4339 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[10]|Q_net  ) );
      defparam \cal1_v__reg[10] .INIT = 0;
      defparam \cal1_v__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[11]  ( .CLK( clkb ), .D( nn4340 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[11]|Q_net  ) );
      defparam \cal1_v__reg[11] .INIT = 0;
      defparam \cal1_v__reg[11] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[12]  ( .CLK( clkb ), .D( nn4341 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[12]|Q_net  ) );
      defparam \cal1_v__reg[12] .INIT = 0;
      defparam \cal1_v__reg[12] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[13]  ( .CLK( clkb ), .D( nn4342 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[13]|Q_net  ) );
      defparam \cal1_v__reg[13] .INIT = 0;
      defparam \cal1_v__reg[13] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[14]  ( .CLK( clkb ), .D( nn4343 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[14]|Q_net  ) );
      defparam \cal1_v__reg[14] .INIT = 0;
      defparam \cal1_v__reg[14] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[15]  ( .CLK( clkb ), .D( nn4344 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[15]|Q_net  ) );
      defparam \cal1_v__reg[15] .INIT = 0;
      defparam \cal1_v__reg[15] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[16]  ( .CLK( clkb ), .D( nn4345 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[16]|Q_net  ) );
      defparam \cal1_v__reg[16] .INIT = 0;
      defparam \cal1_v__reg[16] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[1]  ( .CLK( clkb ), .D( nn4346 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[1]|Q_net  ) );
      defparam \cal1_v__reg[1] .INIT = 0;
      defparam \cal1_v__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[2]  ( .CLK( clkb ), .D( nn4347 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[2]|Q_net  ) );
      defparam \cal1_v__reg[2] .INIT = 0;
      defparam \cal1_v__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[3]  ( .CLK( clkb ), .D( nn4348 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[3]|Q_net  ) );
      defparam \cal1_v__reg[3] .INIT = 0;
      defparam \cal1_v__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[4]  ( .CLK( clkb ), .D( nn4349 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[4]|Q_net  ) );
      defparam \cal1_v__reg[4] .INIT = 0;
      defparam \cal1_v__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[5]  ( .CLK( clkb ), .D( nn4350 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[5]|Q_net  ) );
      defparam \cal1_v__reg[5] .INIT = 0;
      defparam \cal1_v__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[6]  ( .CLK( clkb ), .D( nn4351 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[6]|Q_net  ) );
      defparam \cal1_v__reg[6] .INIT = 0;
      defparam \cal1_v__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[7]  ( .CLK( clkb ), .D( nn4352 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[7]|Q_net  ) );
      defparam \cal1_v__reg[7] .INIT = 0;
      defparam \cal1_v__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[8]  ( .CLK( clkb ), .D( nn4353 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[8]|Q_net  ) );
      defparam \cal1_v__reg[8] .INIT = 0;
      defparam \cal1_v__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_v__reg[9]  ( .CLK( clkb ), .D( nn4354 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_v__reg[9]|Q_net  ) );
      defparam \cal1_v__reg[9] .INIT = 0;
      defparam \cal1_v__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_v__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[0]  ( .CLK( clkb ), .D( nn4355 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[0]|Q_net  ) );
      defparam \cal1_xAddress__reg[0] .INIT = 0;
      defparam \cal1_xAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[10]  ( .CLK( clkb ), .D( nn4380 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[10]|Q_net  ) );
      defparam \cal1_xAddress__reg[10] .INIT = 0;
      defparam \cal1_xAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[1]  ( .CLK( clkb ), .D( nn4381 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[1]|Q_net  ) );
      defparam \cal1_xAddress__reg[1] .INIT = 0;
      defparam \cal1_xAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[2]  ( .CLK( clkb ), .D( nn4382 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[2]|Q_net  ) );
      defparam \cal1_xAddress__reg[2] .INIT = 0;
      defparam \cal1_xAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[3]  ( .CLK( clkb ), .D( nn4383 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[3]|Q_net  ) );
      defparam \cal1_xAddress__reg[3] .INIT = 0;
      defparam \cal1_xAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[4]  ( .CLK( clkb ), .D( nn4384 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[4]|Q_net  ) );
      defparam \cal1_xAddress__reg[4] .INIT = 0;
      defparam \cal1_xAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[5]  ( .CLK( clkb ), .D( nn4385 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[5]|Q_net  ) );
      defparam \cal1_xAddress__reg[5] .INIT = 0;
      defparam \cal1_xAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[6]  ( .CLK( clkb ), .D( nn4386 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[6]|Q_net  ) );
      defparam \cal1_xAddress__reg[6] .INIT = 0;
      defparam \cal1_xAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[7]  ( .CLK( clkb ), .D( nn4387 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[7]|Q_net  ) );
      defparam \cal1_xAddress__reg[7] .INIT = 0;
      defparam \cal1_xAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[8]  ( .CLK( clkb ), .D( nn4388 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[8]|Q_net  ) );
      defparam \cal1_xAddress__reg[8] .INIT = 0;
      defparam \cal1_xAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_xAddress__reg[9]  ( .CLK( clkb ), .D( nn4389 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4283 ), .Q( \cal1_xAddress__reg[9]|Q_net  ) );
      defparam \cal1_xAddress__reg[9] .INIT = 0;
      defparam \cal1_xAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_xAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[0]  ( .CLK( clkb ), .D( nn4390 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[0]|Q_net  ) );
      defparam \cal1_yAddress__reg[0] .INIT = 0;
      defparam \cal1_yAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[10]  ( .CLK( clkb ), .D( nn4415 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[10]|Q_net  ) );
      defparam \cal1_yAddress__reg[10] .INIT = 0;
      defparam \cal1_yAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[1]  ( .CLK( clkb ), .D( nn4416 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[1]|Q_net  ) );
      defparam \cal1_yAddress__reg[1] .INIT = 0;
      defparam \cal1_yAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[2]  ( .CLK( clkb ), .D( nn4417 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[2]|Q_net  ) );
      defparam \cal1_yAddress__reg[2] .INIT = 0;
      defparam \cal1_yAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[3]  ( .CLK( clkb ), .D( nn4418 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[3]|Q_net  ) );
      defparam \cal1_yAddress__reg[3] .INIT = 0;
      defparam \cal1_yAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[4]  ( .CLK( clkb ), .D( nn4419 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[4]|Q_net  ) );
      defparam \cal1_yAddress__reg[4] .INIT = 0;
      defparam \cal1_yAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[5]  ( .CLK( clkb ), .D( nn4420 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[5]|Q_net  ) );
      defparam \cal1_yAddress__reg[5] .INIT = 0;
      defparam \cal1_yAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[6]  ( .CLK( clkb ), .D( nn4421 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[6]|Q_net  ) );
      defparam \cal1_yAddress__reg[6] .INIT = 0;
      defparam \cal1_yAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[7]  ( .CLK( clkb ), .D( nn4422 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[7]|Q_net  ) );
      defparam \cal1_yAddress__reg[7] .INIT = 0;
      defparam \cal1_yAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[8]  ( .CLK( clkb ), .D( nn4423 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[8]|Q_net  ) );
      defparam \cal1_yAddress__reg[8] .INIT = 0;
      defparam \cal1_yAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \cal1_yAddress__reg[9]  ( .CLK( clkb ), .D( nn4424 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn1518 ), .Q( \cal1_yAddress__reg[9]|Q_net  ) );
      defparam \cal1_yAddress__reg[9] .INIT = 0;
      defparam \cal1_yAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \cal1_yAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[0]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[0] .INIT = 0;
      defparam \coefcal1_frameRate__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[1]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[1] .INIT = 0;
      defparam \coefcal1_frameRate__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[2]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[2]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[2] .INIT = 0;
      defparam \coefcal1_frameRate__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[3]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[3] .INIT = 0;
      defparam \coefcal1_frameRate__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[4]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[4] .INIT = 0;
      defparam \coefcal1_frameRate__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[5]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[5]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[5] .INIT = 0;
      defparam \coefcal1_frameRate__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[6]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[6]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[6] .INIT = 0;
      defparam \coefcal1_frameRate__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[7]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[7]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[7] .INIT = 0;
      defparam \coefcal1_frameRate__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_frameRate__reg[8]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_frameRate__reg[8]|Q_net  ) );
      defparam \coefcal1_frameRate__reg[8] .INIT = 0;
      defparam \coefcal1_frameRate__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_frameRate__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM coefcal1_inEn__reg ( .CLK( clka ), .D( nn4425 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_inEn__reg|Q_net  ) );
      defparam coefcal1_inEn__reg.INIT = 0;
      defparam coefcal1_inEn__reg.PLACE_LOCATION = "NONE";
      defparam coefcal1_inEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM coefcal1_work__reg ( .CLK( clka ), .D( nn4527 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_work__reg|Q_net  ) );
      defparam coefcal1_work__reg.INIT = 0;
      defparam coefcal1_work__reg.PLACE_LOCATION = "NONE";
      defparam coefcal1_work__reg.PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[0]|Q_net  ) );
      defparam \coefcal1_working__reg[0] .INIT = 0;
      defparam \coefcal1_working__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[10]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[10]|Q_net  ) );
      defparam \coefcal1_working__reg[10] .INIT = 0;
      defparam \coefcal1_working__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[11]|Q_net  ) );
      defparam \coefcal1_working__reg[11] .INIT = 0;
      defparam \coefcal1_working__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[12]|Q_net  ) );
      defparam \coefcal1_working__reg[12] .INIT = 0;
      defparam \coefcal1_working__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[13]|Q_net  ) );
      defparam \coefcal1_working__reg[13] .INIT = 0;
      defparam \coefcal1_working__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[14]|Q_net  ) );
      defparam \coefcal1_working__reg[14] .INIT = 0;
      defparam \coefcal1_working__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[15]|Q_net  ) );
      defparam \coefcal1_working__reg[15] .INIT = 0;
      defparam \coefcal1_working__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[16]|Q_net  ) );
      defparam \coefcal1_working__reg[16] .INIT = 0;
      defparam \coefcal1_working__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[17]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[17]|Q_net  ) );
      defparam \coefcal1_working__reg[17] .INIT = 0;
      defparam \coefcal1_working__reg[17] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[17] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[18]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[18]|Q_net  ) );
      defparam \coefcal1_working__reg[18] .INIT = 0;
      defparam \coefcal1_working__reg[18] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[18] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[19]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[19]|Q_net  ) );
      defparam \coefcal1_working__reg[19] .INIT = 0;
      defparam \coefcal1_working__reg[19] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[19] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[1]|Q_net  ) );
      defparam \coefcal1_working__reg[1] .INIT = 0;
      defparam \coefcal1_working__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[20]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[20]|Q_net  ) );
      defparam \coefcal1_working__reg[20] .INIT = 0;
      defparam \coefcal1_working__reg[20] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[20] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[21]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[21]|Q_net  ) );
      defparam \coefcal1_working__reg[21] .INIT = 0;
      defparam \coefcal1_working__reg[21] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[21] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[22]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[22]|Q_net  ) );
      defparam \coefcal1_working__reg[22] .INIT = 0;
      defparam \coefcal1_working__reg[22] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[22] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[23]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[23]|Q_net  ) );
      defparam \coefcal1_working__reg[23] .INIT = 0;
      defparam \coefcal1_working__reg[23] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[23] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[24]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[24]|Q_net  ) );
      defparam \coefcal1_working__reg[24] .INIT = 0;
      defparam \coefcal1_working__reg[24] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[24] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[25]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[25]|Q_net  ) );
      defparam \coefcal1_working__reg[25] .INIT = 0;
      defparam \coefcal1_working__reg[25] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[25] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[26]  ( .CLK( clka ), .D( a_dinxy_cen_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[26]|Q_net  ) );
      defparam \coefcal1_working__reg[26] .INIT = 0;
      defparam \coefcal1_working__reg[26] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[26] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[27]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[27]|Q_net  ) );
      defparam \coefcal1_working__reg[27] .INIT = 0;
      defparam \coefcal1_working__reg[27] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[27] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[28]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[28]|Q_net  ) );
      defparam \coefcal1_working__reg[28] .INIT = 0;
      defparam \coefcal1_working__reg[28] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[28] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[29]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[29]|Q_net  ) );
      defparam \coefcal1_working__reg[29] .INIT = 0;
      defparam \coefcal1_working__reg[29] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[29] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[2]|Q_net  ) );
      defparam \coefcal1_working__reg[2] .INIT = 0;
      defparam \coefcal1_working__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[30]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[30]|Q_net  ) );
      defparam \coefcal1_working__reg[30] .INIT = 0;
      defparam \coefcal1_working__reg[30] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[30] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[31]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[31]|Q_net  ) );
      defparam \coefcal1_working__reg[31] .INIT = 0;
      defparam \coefcal1_working__reg[31] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[31] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[32]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[32]|Q_net  ) );
      defparam \coefcal1_working__reg[32] .INIT = 0;
      defparam \coefcal1_working__reg[32] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[32] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[3]|Q_net  ) );
      defparam \coefcal1_working__reg[3] .INIT = 0;
      defparam \coefcal1_working__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[4]|Q_net  ) );
      defparam \coefcal1_working__reg[4] .INIT = 0;
      defparam \coefcal1_working__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[5]|Q_net  ) );
      defparam \coefcal1_working__reg[5] .INIT = 0;
      defparam \coefcal1_working__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[6]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[6]|Q_net  ) );
      defparam \coefcal1_working__reg[6] .INIT = 0;
      defparam \coefcal1_working__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[7]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[7]|Q_net  ) );
      defparam \coefcal1_working__reg[7] .INIT = 0;
      defparam \coefcal1_working__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[8]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[8]|Q_net  ) );
      defparam \coefcal1_working__reg[8] .INIT = 0;
      defparam \coefcal1_working__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_working__reg[9]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_working__reg[9]|Q_net  ) );
      defparam \coefcal1_working__reg[9] .INIT = 0;
      defparam \coefcal1_working__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_working__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[0]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[0] .INIT = 0;
      defparam \coefcal1_xDividend__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[10]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_4|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[10]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[10] .INIT = 0;
      defparam \coefcal1_xDividend__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[11]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_5|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[11]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[11] .INIT = 0;
      defparam \coefcal1_xDividend__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[12]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_6|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[12]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[12] .INIT = 0;
      defparam \coefcal1_xDividend__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[13]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_7|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[13]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[13] .INIT = 0;
      defparam \coefcal1_xDividend__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[14]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_8|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[14]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[14] .INIT = 0;
      defparam \coefcal1_xDividend__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[15]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_9|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[15]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[15] .INIT = 0;
      defparam \coefcal1_xDividend__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[16]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[16]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[16] .INIT = 0;
      defparam \coefcal1_xDividend__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[1]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[1] .INIT = 0;
      defparam \coefcal1_xDividend__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[2]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[2] .INIT = 0;
      defparam \coefcal1_xDividend__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[3]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[3] .INIT = 0;
      defparam \coefcal1_xDividend__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[4]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[4] .INIT = 0;
      defparam \coefcal1_xDividend__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[5]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[5] .INIT = 0;
      defparam \coefcal1_xDividend__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[6]  ( .CLK( clka ), .D( nn4552 ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[6]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[6] .INIT = 0;
      defparam \coefcal1_xDividend__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[7]  ( .CLK( clka ), .D( nn4553 ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[7]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[7] .INIT = 0;
      defparam \coefcal1_xDividend__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[8]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_2|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[8]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[8] .INIT = 0;
      defparam \coefcal1_xDividend__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDividend__reg[9]  ( .CLK( clka ), .D( \coefcal1_u59_XORCI_3|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDividend__reg[9]|Q_net  ) );
      defparam \coefcal1_xDividend__reg[9] .INIT = 0;
      defparam \coefcal1_xDividend__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDividend__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[0]  ( .CLK( clka ), .D( outXRes[0] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[0]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[0] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[10]  ( .CLK( clka ), .D( outXRes[10] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[10]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[10] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[11]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[11] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[12]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[12] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[13]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[13] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[14]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[14] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[15]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[15] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[16]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[16] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[1]  ( .CLK( clka ), .D( outXRes[1] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[1]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[1] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[2]  ( .CLK( clka ), .D( outXRes[2] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[2]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[2] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[3]  ( .CLK( clka ), .D( outXRes[3] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[3]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[3] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[4]  ( .CLK( clka ), .D( outXRes[4] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[4]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[4] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[5]  ( .CLK( clka ), .D( outXRes[5] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[5]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[5] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[6]  ( .CLK( clka ), .D( outXRes[6] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[6]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[6] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[7]  ( .CLK( clka ), .D( outXRes[7] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[7]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[7] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[8]  ( .CLK( clka ), .D( outXRes[8] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[8]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[8] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_xDivisor__reg[9]  ( .CLK( clka ), .D( outXRes[9] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_xDivisor__reg[9]|Q_net  ) );
      defparam \coefcal1_xDivisor__reg[9] .INIT = 0;
      defparam \coefcal1_xDivisor__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_xDivisor__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[0]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[0]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[0] .INIT = 0;
      defparam \coefcal1_yDividend__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[10]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_4|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[10]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[10] .INIT = 0;
      defparam \coefcal1_yDividend__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[11]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_5|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[11]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[11] .INIT = 0;
      defparam \coefcal1_yDividend__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[12]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_6|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[12]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[12] .INIT = 0;
      defparam \coefcal1_yDividend__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[13]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_7|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[13]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[13] .INIT = 0;
      defparam \coefcal1_yDividend__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[14]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_8|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[14]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[14] .INIT = 0;
      defparam \coefcal1_yDividend__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[15]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_9|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[15]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[15] .INIT = 0;
      defparam \coefcal1_yDividend__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[16]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[16]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[16] .INIT = 0;
      defparam \coefcal1_yDividend__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[1]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[1]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[1] .INIT = 0;
      defparam \coefcal1_yDividend__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[2]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[2]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[2] .INIT = 0;
      defparam \coefcal1_yDividend__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[3]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[3]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[3] .INIT = 0;
      defparam \coefcal1_yDividend__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[4]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[4]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[4] .INIT = 0;
      defparam \coefcal1_yDividend__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[5]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[5]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[5] .INIT = 0;
      defparam \coefcal1_yDividend__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[6]  ( .CLK( clka ), .D( nn4604 ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[6]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[6] .INIT = 0;
      defparam \coefcal1_yDividend__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[7]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_1|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[7]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[7] .INIT = 0;
      defparam \coefcal1_yDividend__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[8]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_2|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[8]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[8] .INIT = 0;
      defparam \coefcal1_yDividend__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDividend__reg[9]  ( .CLK( clka ), .D( \coefcal1_u60_XORCI_3|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDividend__reg[9]|Q_net  ) );
      defparam \coefcal1_yDividend__reg[9] .INIT = 0;
      defparam \coefcal1_yDividend__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDividend__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[0]  ( .CLK( clka ), .D( outYRes[0] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[0]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[0] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[0] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[10]  ( .CLK( clka ), .D( outYRes[10] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[10]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[10] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[10] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[10] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[11]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[11]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[11] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[11] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[11] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[12]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[12]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[12] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[12] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[12] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[13]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[13]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[13] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[13] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[13] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[14]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[14]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[14] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[14] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[14] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[15]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[15]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[15] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[15] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[15] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[16]  ( .CLK( clka ), .D( a_acc_en_cal1_u137_mac ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[16]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[16] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[16] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[16] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[1]  ( .CLK( clka ), .D( outYRes[1] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[1]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[1] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[1] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[1] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[2]  ( .CLK( clka ), .D( outYRes[2] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[2]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[2] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[2] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[2] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[3]  ( .CLK( clka ), .D( outYRes[3] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[3]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[3] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[3] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[3] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[4]  ( .CLK( clka ), .D( outYRes[4] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[4]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[4] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[4] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[4] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[5]  ( .CLK( clka ), .D( outYRes[5] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[5]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[5] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[5] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[5] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[6]  ( .CLK( clka ), .D( outYRes[6] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[6]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[6] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[6] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[6] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[7]  ( .CLK( clka ), .D( outYRes[7] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[7]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[7] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[7] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[7] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[8]  ( .CLK( clka ), .D( outYRes[8] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[8]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[8] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[8] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[8] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \coefcal1_yDivisor__reg[9]  ( .CLK( clka ), .D( outYRes[9] ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \coefcal1_yDivisor__reg[9]|Q_net  ) );
      defparam \coefcal1_yDivisor__reg[9] .INIT = 0;
      defparam \coefcal1_yDivisor__reg[9] .PLACE_LOCATION = "NONE";
      defparam \coefcal1_yDivisor__reg[9] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0A_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_0A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_0A_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0A_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0A_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0A_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0A_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_0A_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0A_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0A_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0A_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0B_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_0A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_0A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_0B_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0B_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0B_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0B_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_0B_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_0B_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_0B_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_0B_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_0B_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1A_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_1A_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1A_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1A_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1A_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1A_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_1A_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1A_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1A_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1A_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1B_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_1B_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1B_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1B_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1B_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_1B_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_1B_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_1B_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_1B_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_1B_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3A_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_3A_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3A_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3A_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3A_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3A_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_3A_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3A_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3A_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3A_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3B_aa_reg__reg[0]  ( .CLK( c1r1_clka_fifo1_ram_inst_1A_u_emb18k_0 ), .D( \haa[0]_fifo1_ram_inst_1A_u_emb18k_0  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_3B_aa_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3B_aa_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3B_aa_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3B_aa_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REG_PRIM \fifo1_ram_inst_3B_ab_reg__reg[0]  ( .CLK( clkb ), .D( \cal1_u129_XORCI_10|SUM_net  ), .RST( a_acc_en_cal1_u137_mac ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \fifo1_ram_inst_3B_ab_reg__reg[0]|Q_net  ) );
      defparam \fifo1_ram_inst_3B_ab_reg__reg[0] .INIT = 0;
      defparam \fifo1_ram_inst_3B_ab_reg__reg[0] .PLACE_LOCATION = "NONE";
      defparam \fifo1_ram_inst_3B_ab_reg__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[0]  ( .CLK( clka ), .D( nn4605 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[0]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[0] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[10]  ( .CLK( clka ), .D( nn4728 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[10]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[10] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[11]  ( .CLK( clka ), .D( nn4729 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[11]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[11] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[12]  ( .CLK( clka ), .D( nn4730 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[12]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[12] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[13]  ( .CLK( clka ), .D( nn4731 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[13]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[13] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[14]  ( .CLK( clka ), .D( nn4732 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[14]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[14] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[15]  ( .CLK( clka ), .D( nn4733 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[15]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[15] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[16]  ( .CLK( clka ), .D( nn4734 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[16]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[16] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[16] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[17]  ( .CLK( clka ), .D( nn4735 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[17]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[17] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[17] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[17] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[18]  ( .CLK( clka ), .D( nn4736 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[18]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[18] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[18] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[18] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[19]  ( .CLK( clka ), .D( nn4737 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[19]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[19] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[19] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[19] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[1]  ( .CLK( clka ), .D( nn4738 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[1]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[1] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[20]  ( .CLK( clka ), .D( nn4739 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[20]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[20] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[20] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[20] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[21]  ( .CLK( clka ), .D( nn4740 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[21]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[21] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[21] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[21] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[22]  ( .CLK( clka ), .D( nn4741 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[22]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[22] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[22] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[22] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[23]  ( .CLK( clka ), .D( nn4742 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[23]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[23] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[23] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[23] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[2]  ( .CLK( clka ), .D( nn4743 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[2]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[2] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[3]  ( .CLK( clka ), .D( nn4744 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[3]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[3] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[4]  ( .CLK( clka ), .D( nn4745 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[4]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[4] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[5]  ( .CLK( clka ), .D( nn4746 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[5]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[5] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[6]  ( .CLK( clka ), .D( nn4747 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[6]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[6] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[7]  ( .CLK( clka ), .D( nn4748 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[7]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[7] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[8]  ( .CLK( clka ), .D( nn4749 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[8]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[8] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_dataOut__reg[9]  ( .CLK( clka ), .D( nn4750 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_dataOut__reg[9]|Q_net  ) );
      defparam \inputctrl1_dataOut__reg[9] .INIT = 0;
      defparam \inputctrl1_dataOut__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_dataOut__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_jmp__reg ( .CLK( clka ), .D( nn4751 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4727 ), .Q( \inputctrl1_jmp__reg|Q_net  ) );
      defparam inputctrl1_jmp__reg.INIT = 0;
      defparam inputctrl1_jmp__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_jmp__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[0]  ( .CLK( clka ), .D( nn4752 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[0]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[0] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[10]  ( .CLK( clka ), .D( nn4777 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[10]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[10] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[1]  ( .CLK( clka ), .D( nn4778 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[1]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[1] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[2]  ( .CLK( clka ), .D( nn4779 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[2]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[2] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[3]  ( .CLK( clka ), .D( nn4780 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[3]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[3] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[4]  ( .CLK( clka ), .D( nn4781 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[4]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[4] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[5]  ( .CLK( clka ), .D( nn4782 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[5]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[5] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[6]  ( .CLK( clka ), .D( nn4783 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[6]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[6] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[7]  ( .CLK( clka ), .D( nn4784 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[7]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[7] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[8]  ( .CLK( clka ), .D( nn4785 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[8]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[8] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_ramWrtAddr__reg[9]  ( .CLK( clka ), .D( nn4786 ), .RST( a_acc_en_cal1_u137_mac ), .SET( rst ), .CE( nn4727 ), .Q( \inputctrl1_ramWrtAddr__reg[9]|Q_net  ) );
      defparam \inputctrl1_ramWrtAddr__reg[9] .INIT = 0;
      defparam \inputctrl1_ramWrtAddr__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_ramWrtAddr__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_ramWrtEn__reg ( .CLK( clka ), .D( nn4787 ), .RST( rst ), .SET( a_acc_en_cal1_u137_mac ), .CE( a_dinxy_cen_cal1_u137_mac ), .Q( \inputctrl1_ramWrtEn__reg|Q_net  ) );
      defparam inputctrl1_ramWrtEn__reg.INIT = 0;
      defparam inputctrl1_ramWrtEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_ramWrtEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[0]  ( .CLK( clka ), .D( nn4788 ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[0]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[0] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_10|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[10]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[10] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_1|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[1]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[1] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_2|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[2]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[2] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_3|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[3]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[3] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_4|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[4]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[4] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_5|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[5]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[5] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_6|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[6]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[6] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_7|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[7]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[7] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_8|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[8]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[8] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xAddress__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u110_XORCI_9|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xAddress__reg[9]|Q_net  ) );
      defparam \inputctrl1_xAddress__reg[9] .INIT = 0;
      defparam \inputctrl1_xAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[0]  ( .CLK( clka ), .D( nn4816 ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[0]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[0] .INIT = 0;
      defparam \inputctrl1_xCal__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_10|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[10]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[10] .INIT = 0;
      defparam \inputctrl1_xCal__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[11]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_11|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[11]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[11] .INIT = 0;
      defparam \inputctrl1_xCal__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[12]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_12|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[12]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[12] .INIT = 0;
      defparam \inputctrl1_xCal__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[13]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_13|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[13]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[13] .INIT = 0;
      defparam \inputctrl1_xCal__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[14]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_14|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[14]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[14] .INIT = 0;
      defparam \inputctrl1_xCal__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[15]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_15|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[15]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[15] .INIT = 0;
      defparam \inputctrl1_xCal__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[16]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_16|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[16]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[16] .INIT = 0;
      defparam \inputctrl1_xCal__reg[16] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_1|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[1]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[1] .INIT = 0;
      defparam \inputctrl1_xCal__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_2|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[2]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[2] .INIT = 0;
      defparam \inputctrl1_xCal__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_3|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[3]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[3] .INIT = 0;
      defparam \inputctrl1_xCal__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_4|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[4]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[4] .INIT = 0;
      defparam \inputctrl1_xCal__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_5|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[5]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[5] .INIT = 0;
      defparam \inputctrl1_xCal__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_6|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[6]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[6] .INIT = 0;
      defparam \inputctrl1_xCal__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_7|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[7]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[7] .INIT = 0;
      defparam \inputctrl1_xCal__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_8|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[8]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[8] .INIT = 0;
      defparam \inputctrl1_xCal__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_xCal__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u108_XORCI_9|SUM_net  ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4817 ), .Q( \inputctrl1_xCal__reg[9]|Q_net  ) );
      defparam \inputctrl1_xCal__reg[9] .INIT = 0;
      defparam \inputctrl1_xCal__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_xCal__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_xPreEn__reg ( .CLK( clka ), .D( nn4612 ), .RST( nn4789 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4790 ), .Q( \inputctrl1_xPreEn__reg|Q_net  ) );
      defparam inputctrl1_xPreEn__reg.INIT = 0;
      defparam inputctrl1_xPreEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_xPreEn__reg.PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[0]  ( .CLK( clka ), .D( nn4854 ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[0]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[0] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_10|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[10]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[10] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_1|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[1]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[1] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_2|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[2]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[2] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_3|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[3]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[3] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_4|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[4]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[4] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_5|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[5]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[5] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_6|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[6]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[6] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_7|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[7]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[7] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_8|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[8]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[8] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yAddress__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u111_XORCI_9|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yAddress__reg[9]|Q_net  ) );
      defparam \inputctrl1_yAddress__reg[9] .INIT = 0;
      defparam \inputctrl1_yAddress__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yAddress__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[0]  ( .CLK( clka ), .D( nn4881 ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[0]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[0] .INIT = 0;
      defparam \inputctrl1_yCal__reg[0] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[0] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[10]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_10|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[10]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[10] .INIT = 0;
      defparam \inputctrl1_yCal__reg[10] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[10] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[11]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_11|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[11]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[11] .INIT = 0;
      defparam \inputctrl1_yCal__reg[11] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[11] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[12]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_12|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[12]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[12] .INIT = 0;
      defparam \inputctrl1_yCal__reg[12] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[12] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[13]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_13|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[13]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[13] .INIT = 0;
      defparam \inputctrl1_yCal__reg[13] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[13] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[14]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_14|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[14]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[14] .INIT = 0;
      defparam \inputctrl1_yCal__reg[14] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[14] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[15]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_15|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[15]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[15] .INIT = 0;
      defparam \inputctrl1_yCal__reg[15] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[15] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[16]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_16|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[16]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[16] .INIT = 0;
      defparam \inputctrl1_yCal__reg[16] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[16] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[1]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_1|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[1]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[1] .INIT = 0;
      defparam \inputctrl1_yCal__reg[1] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[1] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[2]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_2|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[2]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[2] .INIT = 0;
      defparam \inputctrl1_yCal__reg[2] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[2] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[3]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_3|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[3]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[3] .INIT = 0;
      defparam \inputctrl1_yCal__reg[3] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[3] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[4]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_4|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[4]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[4] .INIT = 0;
      defparam \inputctrl1_yCal__reg[4] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[4] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[5]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_5|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[5]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[5] .INIT = 0;
      defparam \inputctrl1_yCal__reg[5] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[5] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[6]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_6|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[6]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[6] .INIT = 0;
      defparam \inputctrl1_yCal__reg[6] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[6] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[7]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_7|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[7]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[7] .INIT = 0;
      defparam \inputctrl1_yCal__reg[7] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[7] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[8]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_8|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[8]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[8] .INIT = 0;
      defparam \inputctrl1_yCal__reg[8] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[8] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM \inputctrl1_yCal__reg[9]  ( .CLK( clka ), .D( \inputctrl1_u109_XORCI_9|SUM_net  ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( nn4882 ), .Q( \inputctrl1_yCal__reg[9]|Q_net  ) );
      defparam \inputctrl1_yCal__reg[9] .INIT = 0;
      defparam \inputctrl1_yCal__reg[9] .PLACE_LOCATION = "NONE";
      defparam \inputctrl1_yCal__reg[9] .PCK_LOCATION = "NONE";
    CS_REGA_PRIM inputctrl1_yPreEn__reg ( .CLK( clka ), .D( nn4645 ), .RST( nn4855 ), .SET( a_acc_en_cal1_u137_mac ), .CE( iHsyn ), .Q( \inputctrl1_yPreEn__reg|Q_net  ) );
      defparam inputctrl1_yPreEn__reg.INIT = 0;
      defparam inputctrl1_yPreEn__reg.PLACE_LOCATION = "NONE";
      defparam inputctrl1_yPreEn__reg.PCK_LOCATION = "NONE";

endmodule


