.box 1 scaler_ipc_adder_17 35 18
.input 1 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16]
.output 1 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] CO
.delay 1
-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	1200	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1300	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1400	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1500	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1600	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1700	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1800	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 2 scaler_ipc_adder_11 23 12
.input 2 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10]
.output 2 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] CO
.delay 2
-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	
1000	900	800	700	600	500	400	300	200	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	
1100	1000	900	800	700	600	500	400	300	200	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	
1200	1100	1000	900	800	700	600	500	400	300	200	1200	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 3 scaler_ipc_adder_7 15 8
.input 3 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6]
.output 3 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] CO
.delay 3
-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	
200	-	-	-	-	-	-	200	200	100	-	-	-	-	-	
300	200	-	-	-	-	-	300	300	200	100	-	-	-	-	
400	300	200	-	-	-	-	400	400	300	200	100	-	-	-	
500	400	300	200	-	-	-	500	500	400	300	200	100	-	-	
600	500	400	300	200	-	-	600	600	500	400	300	200	100	-	
700	600	500	400	300	200	-	700	700	600	500	400	300	200	100	
800	700	600	500	400	300	200	800	800	700	600	500	400	300	200	


.box 4 scaler_ipc_adder_9 19 10
.input 4 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8]
.output 4 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] CO
.delay 4
-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	
600	500	400	300	200	-	-	-	-	600	600	500	400	300	200	100	-	-	-	
700	600	500	400	300	200	-	-	-	700	700	600	500	400	300	200	100	-	-	
800	700	600	500	400	300	200	-	-	800	800	700	600	500	400	300	200	100	-	
900	800	700	600	500	400	300	200	-	900	900	800	700	600	500	400	300	200	100	
1000	900	800	700	600	500	400	300	200	1000	1000	900	800	700	600	500	400	300	200	


.box 5 scaler_ipc_adder_10 21 11
.input 5 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9]
.output 5 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] CO
.delay 5
-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	
800	700	600	500	400	300	200	-	-	-	800	800	700	600	500	400	300	200	100	-	-	
900	800	700	600	500	400	300	200	-	-	900	900	800	700	600	500	400	300	200	100	-	
1000	900	800	700	600	500	400	300	200	-	1000	1000	900	800	700	600	500	400	300	200	100	
1100	1000	900	800	700	600	500	400	300	200	1100	1100	1000	900	800	700	600	500	400	300	200	


.box 6 scaler_ipc_adder_12 25 13
.input 6 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11]
.output 6 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] CO
.delay 6
-	-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	1200	1200	1100	1000	900	800	700	600	500	400	300	200	100	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	1300	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 7 scaler_ipc_adder_18 37 19
.input 7 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CA[17] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16] DX[17]
.output 7 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] SUM[17] CO
.delay 7
-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	1200	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	1300	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1400	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1500	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1600	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1700	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1800	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1900	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 8 scaler_ipc_adder_8 17 9
.input 8 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7]
.output 8 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] CO
.delay 8
-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	
400	300	200	-	-	-	-	-	400	400	300	200	100	-	-	-	-	
500	400	300	200	-	-	-	-	500	500	400	300	200	100	-	-	-	
600	500	400	300	200	-	-	-	600	600	500	400	300	200	100	-	-	
700	600	500	400	300	200	-	-	700	700	600	500	400	300	200	100	-	
800	700	600	500	400	300	200	-	800	800	700	600	500	400	300	200	100	
900	800	700	600	500	400	300	200	900	900	800	700	600	500	400	300	200	


.box 9 scaler_ipc_adder_14 29 15
.input 9 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13]
.output 9 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] CO
.delay 9
-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	1200	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	1300	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	1400	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	1500	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


.box 10 scaler_ipc_adder_34 69 35
.input 10 CA[0] CA[1] CA[2] CA[3] CA[4] CA[5] CA[6] CA[7] CA[8] CA[9] CA[10] CA[11] CA[12] CA[13] CA[14] CA[15] CA[16] CA[17] CA[18] CA[19] CA[20] CA[21] CA[22] CA[23] CA[24] CA[25] CA[26] CA[27] CA[28] CA[29] CA[30] CA[31] CA[32] CA[33] CI DX[0] DX[1] DX[2] DX[3] DX[4] DX[5] DX[6] DX[7] DX[8] DX[9] DX[10] DX[11] DX[12] DX[13] DX[14] DX[15] DX[16] DX[17] DX[18] DX[19] DX[20] DX[21] DX[22] DX[23] DX[24] DX[25] DX[26] DX[27] DX[28] DX[29] DX[30] DX[31] DX[32] DX[33]
.output 10 SUM[0] SUM[1] SUM[2] SUM[3] SUM[4] SUM[5] SUM[6] SUM[7] SUM[8] SUM[9] SUM[10] SUM[11] SUM[12] SUM[13] SUM[14] SUM[15] SUM[16] SUM[17] SUM[18] SUM[19] SUM[20] SUM[21] SUM[22] SUM[23] SUM[24] SUM[25] SUM[26] SUM[27] SUM[28] SUM[29] SUM[30] SUM[31] SUM[32] SUM[33] CO
.delay 10
-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	100	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	200	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	300	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	400	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	500	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	600	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	700	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	800	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	900	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1000	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1100	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1200	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1300	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1400	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1500	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1600	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1700	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1800	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	1900	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	-	2000	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	-	
2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	-	2100	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	-	
2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	-	2200	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	-	
2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	-	2300	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	-	
2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	-	2400	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	-	
2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	-	2500	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	-	
2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	-	2600	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	-	
2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	-	2700	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	-	
2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	-	2800	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	-	
2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	-	2900	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	-	
3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	-	3000	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	-	
3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	-	3100	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	-	
3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	-	3200	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	-	
3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	-	3300	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	-	
3400	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	-	3400	3400	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	100	
3500	3400	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	3500	3500	3400	3300	3200	3100	3000	2900	2800	2700	2600	2500	2400	2300	2200	2100	2000	1900	1800	1700	1600	1500	1400	1300	1200	1100	1000	900	800	700	600	500	400	300	200	


