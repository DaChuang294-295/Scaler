library verilog;
use verilog.vl_types.all;
entity DELAY_BUF is
    port(
        \in\            : in     vl_logic;
        \out\           : out    vl_logic
    );
end DELAY_BUF;
